
module alu ( a, b, ALUCtrl, out, zero_signal );
  input [0:31] a;
  input [0:31] b;
  input [0:3] ALUCtrl;
  output [0:31] out;
  output zero_signal;
  wire   n24, n620, n716, n853, n890, n949, n1323, n1386, n1671, n3662,
         net240761, net240762, net240767, net240772, net240774, net240775,
         net240782, net240783, net240784, net240812, net240813, net240814,
         net240839, net240852, net240910, net240912, net240913, net240915,
         net240917, net240927, net240928, net240941, net240951, net240952,
         net240961, net240975, net240978, net240980, net240981, net240982,
         net240985, net240986, net240988, net240989, net240990, net240991,
         net240992, net240994, net240995, net240996, net240997, net241012,
         net241013, net241014, net241021, net241026, net241030, net241031,
         net241032, net241036, net241038, net241039, net241040, net241042,
         net241044, net241045, net241047, net241048, net241050, net241052,
         net241053, net241061, net241062, net241064, net241065, net241069,
         net241072, net241073, net241276, net241491, net241492, net241493,
         net241503, net241542, net241554, net241561, net241562, net241563,
         net241565, net241566, net241567, net241568, net241579, net241581,
         net241596, net241597, net241598, net241599, net241600, net241613,
         net241625, net241628, net241746, net241749, net241751, net241754,
         net241756, net241757, net241758, net241760, net241767, net241770,
         net241771, net241773, net241814, net241817, net241821, net241824,
         net241826, net241827, net241828, net241829, net241830, net241831,
         net241832, net242066, net242067, net242074, net242076, net242079,
         net242080, net242095, net242097, net242098, net242099, net242102,
         net242103, net242110, net242151, net242153, net242309, net242310,
         net242311, net242313, net242315, net242316, net242319, net242322,
         net242324, net242361, net242366, net242367, net242378, net242379,
         net242385, net242402, net242580, net242581, net242594, net242595,
         net242597, net242602, net242611, net242655, net242658, net242659,
         net242666, net242672, net242674, net242810, net242811, net242812,
         net242813, net242817, net242819, net242821, net242823, net242824,
         net242877, net242878, net242879, net242882, net242883, net242885,
         net242894, net242896, net242898, net242899, net242900, net242904,
         net242906, net242907, net242908, net242909, net242910, net242911,
         net242916, net242917, net243066, net243078, net243079, net243080,
         net243081, net243093, net243094, net243096, net243098, net243099,
         net243106, net243118, net243119, net243159, net243164, net243166,
         net243167, net243168, net243171, net243172, net243175, net243176,
         net243177, net243179, net243182, net243184, net243187, net243261,
         net243268, net243270, net243271, net243275, net243277, net243278,
         net243279, net243281, net243283, net243284, net243286, net243288,
         net243289, net243291, net243292, net243293, net243294, net243296,
         net243298, net243299, net243310, net243311, net243356, net243367,
         net243368, net243371, net243374, net243376, net243395, net243396,
         net243398, net243399, net243400, net243403, net243404, net243405,
         net243406, net243422, net243423, net243433, net243439, net243578,
         net243582, net243584, net243587, net243625, net243628, net243630,
         net243634, net243637, net243639, net243645, net243723, net243725,
         net243727, net243731, net243733, net243734, net243740, net243741,
         net243743, net243747, net243754, net243755, net243757, net243759,
         net243760, net243761, net243763, net243765, net243769, net243770,
         net243771, net243774, net243775, net243778, net243781, net243785,
         net243790, net243791, net243844, net243866, net243868, net243991,
         net243999, net244001, net244005, net244006, net244008, net244055,
         net244056, net244062, net244063, net244064, net244072, net244073,
         net244074, net244075, net244076, net244078, net244136, net244143,
         net244144, net244145, net244156, net244173, net244177, net244178,
         net244180, net244181, net244239, net244243, net244244, net244256,
         net244257, net244258, net244260, net244262, net244271, net244272,
         net244278, net244281, net244283, net244284, net244285, net244287,
         net244288, net244368, net244369, net244370, net244371, net244373,
         net244374, net244384, net244442, net244457, net244522, net244523,
         net244528, net244529, net244535, net244537, net244540, net244541,
         net244543, net244545, net244546, net244554, net244567, net244568,
         net244627, net244655, net244659, net244665, net244666, net244669,
         net244674, net244679, net244681, net244682, net244683, net244686,
         net244688, net244689, net244690, net244701, net244702, net244704,
         net244808, net244841, net244862, net244867, net244872, net244873,
         net244874, net244875, net244933, net245029, net245052, net245207,
         net245209, net245249, net245250, net245266, net245268, net245313,
         net245317, net245318, net245348, net245349, net245359, net245369,
         net245387, net245388, net245389, net245393, net245422, net245429,
         net245459, net245465, net245474, net245501, net245523, net245524,
         net245525, net245541, net245546, net245611, net245614, net245615,
         net245617, net245621, net245672, net245673, net245674, net245675,
         net245697, net245698, net245700, net245702, net245703, net245711,
         net245722, net245724, net245731, net245732, net245737, net245738,
         net245739, net245740, net245741, net245742, net245752, net245760,
         net245761, net245762, net245764, net245765, net245768, net245774,
         net245775, net245782, net245783, net245785, net245786, net245794,
         net245799, net245800, net245801, net245802, net245803, net245804,
         net245805, net245806, net245808, net245809, net245810, net245888,
         net245906, net245907, net245909, net245910, net245911, net245918,
         net245919, net245920, net245921, net245959, net245960, net245962,
         net245963, net245981, net245984, net245985, net245988, net245989,
         net245991, net245992, net246003, net246013, net246014, net246016,
         net246017, net246031, net246034, net246068, net246070, net246071,
         net246072, net246073, net246074, net246075, net246076, net246077,
         net246082, net246086, net246089, net246091, net246096, net246100,
         net246105, net246106, net246107, net246116, net246117, net246118,
         net246120, net246127, net246129, net246130, net246131, net246132,
         net246133, net246135, net246172, net246176, net246177, net246179,
         net246181, net246186, net246188, net246190, net246198, net246204,
         net246205, net246235, net246238, net246239, net246244, net246250,
         net246254, net246272, net246273, net246274, net246287, net246288,
         net246289, net246327, net246332, net246342, net246345, net246346,
         net246348, net246349, net246353, net246381, net246382, net246384,
         net246385, net246386, net246387, net246389, net246392, net246393,
         net246395, net246397, net246401, net246402, net246403, net246407,
         net246431, net246432, net246433, net246434, net246443, net246445,
         net246446, net246447, net246448, net246450, net246463, net246466,
         net246470, net246475, net246481, net246482, net246483, net246497,
         net246506, net246509, net246511, net246513, net246514, net246515,
         net246525, net246530, net246534, net246535, net246536, net246539,
         net246542, net246545, net246552, net246557, net246558, net246564,
         net246566, net246569, net246570, net246576, net246577, net246578,
         net246579, net246589, net246750, net246756, net246754, net246764,
         net246762, net246760, net246770, net246768, net246766, net246776,
         net246772, net246782, net246792, net246790, net246788, net246786,
         net246804, net246812, net246832, net246836, net246844, net246850,
         net246862, net246868, net246876, net246874, net246888, net246886,
         net246882, net246880, net246878, net246908, net246904, net246902,
         net246920, net246918, net246916, net246932, net246930, net246926,
         net246924, net246958, net246956, net246966, net246962, net246960,
         net246970, net247002, net247044, net247043, net247049, net247048,
         net247060, net247059, net247083, net247082, net247168, net247167,
         net247473, net247540, net247545, net247549, net247630, net247632,
         net247660, net247659, net247658, net247741, net247752, net247751,
         net247762, net247778, net247821, net247820, net247817, net247815,
         net247809, net247808, net247807, net247804, net247843, net247847,
         net247881, net248031, net248030, net248029, net248040, net248038,
         net248078, net248083, net248207, net248350, net248354, net248353,
         net248371, net248379, net248395, net248403, net248433, net248432,
         net248442, net248444, net248449, net248509, net248511, net248517,
         net248516, net248549, net248615, net248620, net248639, net248651,
         net248693, net248717, net248742, net248749, net248775, net248776,
         net248780, net248788, net248893, net248913, net248925, net248960,
         net248987, net248988, net249059, net249076, net249104, net249128,
         net249130, net249142, net249177, net249183, net249187, net249194,
         net249225, net249231, net249298, net249316, net249328, net249335,
         net249352, net249197, net244695, net244668, net244565, net246251,
         net243863, net243776, net242839, net242835, net246838, net244687,
         net244684, net241614, net241607, net246778, net241582, net241573,
         net240983, net240960, net240958, net240956, net243375, net243373,
         net243185, net242314, net240925, net240916, net246516, net246510,
         net246468, net243290, net243101, net243100, net243082, net242604,
         net242818, net244465, net244274, net244273, net242068, net241772,
         net241020, net240930, net240929, net247211, net247164, net244671,
         net244667, net244555, net244553, net249297, net243108, net242830,
         net242826, net247173, net246551, net243636, net243635, net243583,
         net246008, net246007, net246005, net246559, net247667, net246582,
         net246394, net246390, net246361, net246359, net246237, net248923,
         net246199, net243990, net243989, net243728, net244077, net245896,
         net245895, net245893, net245892, net245756, net243652, net243580,
         net243401, net243301, net243300, net243297, net242321, net242305,
         net242304, net242303, net246526, net246523, net248703, net243181,
         net247223, net243875, net243777, net243729, net243726, net248389,
         net247491, net245734, net245616, net244698, net244697, net244696,
         net244692, net244685, net241010, net248477, net243651, net243579,
         net243392, net243391, net243378, net243308, net243307, net243295,
         net243285, net241024, net241023, net246081, net246080, net245993,
         net245766, net245759, net246269, net248217, net248216, net246281,
         net246277, net246275, net246248, net246243, net246236, net249278,
         net249044, net249043, net248695, net241033, net241029, net240999,
         net240949, net240939, net240937, net240936, net240924, net242837,
         net247563, net244066, net243780, net241070, net241063, net245730,
         net245613, net245612, net244564, net244563, net244562, net244561,
         net244560, net244559, net244558, net244557, net246518, net246502,
         net246485, net246452, net248692, net241587, net241071, net241022,
         net241018, net241011, net241009, net241006, net248132, net245897,
         net248551, net247924, net244379, net244270, net244154, net244152,
         net244151, net244150, net240966, net240962, net240954, net240953,
         net240944, net240934, net240933, net240932, net240931, net244067,
         net243995, net243988, net246974, net240918, net240763, net246114,
         net246113, net246002, net249302, net248623, net246206, net246000,
         net246437, net246400, net246396, net246581, net245690, net245689,
         net245686, net245679, net246006, net247544, net244372, net244289,
         net244146, net249331, net245680, net245678, net245677, net244694,
         net246262, net246261, net246260, net246258, net246201, net246200,
         net246111, net246109, net246004, net241007, net241005, net241003,
         net241002, net248357, net245956, net245955, net245954, net245953,
         net245952, net245773, net245757, net248400, net247919, net247918,
         net247917, net247916, net243105, net243104, net242901, net242832,
         net242829, net242828, net242827, net242825, net242822, net243631,
         net243362, net243313, net243186, net249149, net246910, net246541,
         net246540, net249300, net248867, net248865, net248612, net245890,
         net245751, net245750, net245745, net245744, net245691, net243998,
         net243997, net243996, net243860, net243784, net243782, net243408,
         net242323, net241612, net249274, net248800, net246856, net246110,
         net246108, net245998, net245902, net245901, net245899, net245898,
         net244378, net244269, net244263, net244163, net244161, net244160,
         net244153, net243994, net246568, net246561, net246560, net246544,
         net246543, net246538, net246537, net242072, net242071, net241608,
         net248443, net247850, net243874, net243865, net243862, net243861,
         net243789, net243788, net243787, net243779, net243407, net248571,
         net246491, net246488, net243377, net243370, net243369, net243361,
         net243315, net243314, net243180, net243121, net243114, net243113,
         net243111, net243110, net242838, net242836, net242833, net242831,
         net248778, net248777, net247915, net242891, net242884, net242834,
         net242673, net242669, net242668, net242613, net242612, net242610,
         net242609, net242608, net242607, net242606, net242605, net242603,
         net248472, net245758, net245755, net245754, net245753, net245696,
         net245694, net245688, net245687, net245683, net245681, net245676,
         net244155, net243993, net243749, net243746, net243745, net241595,
         net241594, net241593, net247928, net247927, net247926, net244466,
         net244387, net244386, net244385, net244383, net244382, net244381,
         net244380, net244275, net246439, net246438, net246388, net247619,
         net246436, net246365, net246364, net246363, net246362, net246360,
         net246358, net246357, net246247, net246246, net246242, net246241,
         net249292, net242667, net242383, net242382, net242377, net242376,
         net242375, net242368, net242325, net242320, net242302, net242101,
         net242100, net241004, net241001, net241000, net240965, net240964,
         net240963, net247186, net246550, net246549, net246521, net246520,
         net245997, net245994, net245958, net245957, net245905, net245904,
         net247797, net247795, net246522, net246517, net246487, net246486,
         net246484, net246480, net246479, net246478, net246477, net246476,
         net246467, net246399, net246398, net247912, net242077, net242070,
         net242069, net241616, net241615, net241611, net241610, net241609,
         net241606, net241589, net241588, net241586, net241068, net241067,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868;

  AOI21_X4 U601 ( .B1(net246960), .B2(a[7]), .A(n24), .ZN(n853) );
  AOI21_X4 U908 ( .B1(net246960), .B2(a[3]), .A(n24), .ZN(n1386) );
  AOI21_X4 U912 ( .B1(net246960), .B2(a[4]), .A(n24), .ZN(n949) );
  AOI21_X4 U2938 ( .B1(net246960), .B2(a[0]), .A(n24), .ZN(n1323) );
  NOR2_X4 U3191 ( .A1(n4566), .A2(net246956), .ZN(n1671) );
  NOR2_X4 U3220 ( .A1(b[29]), .A2(net248516), .ZN(n716) );
  NOR2_X4 U3226 ( .A1(b[27]), .A2(net246878), .ZN(n890) );
  INV_X4 U3848 ( .A(n1671), .ZN(n620) );
  INV_X2 U3878 ( .A(net245920), .ZN(n4338) );
  INV_X4 U3879 ( .A(net245810), .ZN(net245809) );
  NAND2_X2 U3880 ( .A1(n4504), .A2(n4505), .ZN(n5937) );
  NAND2_X1 U3881 ( .A1(net242098), .A2(net241613), .ZN(n3847) );
  NAND2_X2 U3882 ( .A1(n3845), .A2(n3846), .ZN(n3848) );
  NAND2_X2 U3883 ( .A1(n3847), .A2(n3848), .ZN(n7860) );
  INV_X2 U3884 ( .A(net242098), .ZN(n3845) );
  INV_X1 U3885 ( .A(net241613), .ZN(n3846) );
  NAND2_X4 U3886 ( .A1(a[2]), .A2(b[31]), .ZN(n8352) );
  NAND2_X4 U3887 ( .A1(a[3]), .A2(b[31]), .ZN(n8195) );
  NAND2_X4 U3888 ( .A1(a[4]), .A2(b[31]), .ZN(n8197) );
  NAND2_X4 U3889 ( .A1(a[5]), .A2(b[31]), .ZN(n7719) );
  NAND2_X4 U3890 ( .A1(a[6]), .A2(b[31]), .ZN(n7721) );
  NAND2_X4 U3891 ( .A1(a[7]), .A2(b[31]), .ZN(n7315) );
  NAND2_X4 U3892 ( .A1(a[9]), .A2(b[31]), .ZN(n6969) );
  INV_X8 U3893 ( .A(net241012), .ZN(n3888) );
  NAND2_X1 U3894 ( .A1(net247778), .A2(net246327), .ZN(n3849) );
  XNOR2_X2 U3895 ( .A(n3851), .B(n3850), .ZN(n7154) );
  INV_X32 U3896 ( .A(n7147), .ZN(n3850) );
  XNOR2_X2 U3897 ( .A(n7145), .B(n7144), .ZN(n3851) );
  INV_X1 U3898 ( .A(n6746), .ZN(n6670) );
  NAND2_X1 U3899 ( .A1(n8070), .A2(n7702), .ZN(n8073) );
  OAI21_X2 U3900 ( .B1(n6958), .B2(n7089), .A(n7094), .ZN(n7098) );
  INV_X4 U3901 ( .A(n4042), .ZN(net241610) );
  AOI21_X4 U3902 ( .B1(net244535), .B2(n6032), .A(net244537), .ZN(n6034) );
  INV_X4 U3903 ( .A(n6822), .ZN(n4480) );
  NAND2_X4 U3904 ( .A1(n5030), .A2(n5029), .ZN(n5037) );
  INV_X4 U3905 ( .A(net244275), .ZN(net247926) );
  NAND2_X4 U3906 ( .A1(n4495), .A2(net247815), .ZN(n5284) );
  NAND2_X4 U3907 ( .A1(net246272), .A2(net246274), .ZN(n4741) );
  INV_X4 U3908 ( .A(n4015), .ZN(n3852) );
  INV_X2 U3909 ( .A(n4015), .ZN(net246242) );
  INV_X8 U3910 ( .A(n7598), .ZN(n7370) );
  INV_X2 U3911 ( .A(net240958), .ZN(net240983) );
  OAI22_X2 U3912 ( .A1(n3897), .A2(n7459), .B1(n7459), .B2(n7458), .ZN(n7461)
         );
  INV_X2 U3913 ( .A(net241073), .ZN(net241276) );
  INV_X2 U3914 ( .A(n4353), .ZN(n6939) );
  NAND2_X2 U3915 ( .A1(n6726), .A2(net243578), .ZN(n6730) );
  AOI211_X1 U3916 ( .C1(n7823), .C2(net246974), .A(n7822), .B(n4267), .ZN(
        n7854) );
  NAND2_X4 U3917 ( .A1(net241022), .A2(net241040), .ZN(net241036) );
  NAND2_X4 U3918 ( .A1(net241616), .A2(net241615), .ZN(net241067) );
  INV_X2 U3919 ( .A(net241616), .ZN(net242069) );
  NAND2_X2 U3920 ( .A1(net249335), .A2(net246089), .ZN(n3855) );
  NAND2_X4 U3921 ( .A1(n3853), .A2(n3854), .ZN(n3856) );
  NAND2_X2 U3922 ( .A1(n3855), .A2(n3856), .ZN(n4878) );
  INV_X4 U3923 ( .A(net249335), .ZN(n3853) );
  INV_X2 U3924 ( .A(net246089), .ZN(n3854) );
  NAND2_X4 U3925 ( .A1(b[23]), .A2(a[28]), .ZN(net246089) );
  NAND2_X1 U3926 ( .A1(n4698), .A2(n4766), .ZN(n4692) );
  AOI21_X2 U3927 ( .B1(net248207), .B2(net245750), .A(net245751), .ZN(n4206)
         );
  INV_X2 U3928 ( .A(net242101), .ZN(n3895) );
  INV_X4 U3929 ( .A(net247563), .ZN(n3918) );
  NAND2_X4 U3930 ( .A1(n3869), .A2(n3870), .ZN(n3872) );
  NAND2_X2 U3931 ( .A1(n4794), .A2(n4793), .ZN(n3859) );
  NAND2_X4 U3932 ( .A1(n3857), .A2(n3858), .ZN(n3860) );
  NAND2_X4 U3933 ( .A1(n3859), .A2(n3860), .ZN(net246129) );
  INV_X4 U3934 ( .A(n4794), .ZN(n3857) );
  INV_X2 U3935 ( .A(n4793), .ZN(n3858) );
  NAND2_X2 U3936 ( .A1(net243391), .A2(net243392), .ZN(n3863) );
  NAND2_X4 U3937 ( .A1(n3861), .A2(n3862), .ZN(n3864) );
  NAND2_X4 U3938 ( .A1(n3863), .A2(n3864), .ZN(net243308) );
  INV_X4 U3939 ( .A(net243391), .ZN(n3861) );
  INV_X4 U3940 ( .A(net243392), .ZN(n3862) );
  NAND2_X2 U3941 ( .A1(n4329), .A2(net245892), .ZN(n3867) );
  NAND2_X4 U3942 ( .A1(n3865), .A2(n3866), .ZN(n3868) );
  NAND2_X4 U3943 ( .A1(n3867), .A2(n3868), .ZN(net245756) );
  INV_X4 U3944 ( .A(n4329), .ZN(n3865) );
  INV_X4 U3945 ( .A(net245892), .ZN(n3866) );
  INV_X8 U3946 ( .A(net243308), .ZN(net243377) );
  NAND2_X4 U3947 ( .A1(net245758), .A2(net245756), .ZN(net245753) );
  NAND2_X1 U3948 ( .A1(n4176), .A2(net243181), .ZN(n3871) );
  NAND2_X2 U3949 ( .A1(n3871), .A2(n3872), .ZN(net243369) );
  INV_X4 U3950 ( .A(n4176), .ZN(n3869) );
  INV_X1 U3951 ( .A(net243181), .ZN(n3870) );
  NAND2_X2 U3952 ( .A1(net241022), .A2(n4278), .ZN(n3875) );
  NAND2_X4 U3953 ( .A1(n3873), .A2(n3874), .ZN(n3876) );
  NAND2_X4 U3954 ( .A1(n3875), .A2(n3876), .ZN(net248692) );
  INV_X2 U3955 ( .A(net241022), .ZN(n3873) );
  INV_X4 U3956 ( .A(n4278), .ZN(n3874) );
  NOR2_X4 U3957 ( .A1(net248692), .A2(net241009), .ZN(net241005) );
  NAND2_X4 U3958 ( .A1(net241009), .A2(net248692), .ZN(net241007) );
  NAND2_X1 U3959 ( .A1(n7816), .A2(n7815), .ZN(n7863) );
  XNOR2_X2 U3960 ( .A(n4722), .B(n4764), .ZN(n4085) );
  NAND2_X4 U3961 ( .A1(n6081), .A2(n6080), .ZN(n5906) );
  INV_X4 U3962 ( .A(n7862), .ZN(n7641) );
  NAND2_X4 U3963 ( .A1(n4998), .A2(n4997), .ZN(n5094) );
  NOR2_X4 U3964 ( .A1(n6210), .A2(n6209), .ZN(n6213) );
  NOR3_X4 U3965 ( .A1(n4462), .A2(n7462), .A3(n7461), .ZN(n7467) );
  INV_X2 U3966 ( .A(n4067), .ZN(n4061) );
  NAND2_X4 U3967 ( .A1(n3994), .A2(n8772), .ZN(net240941) );
  NAND2_X4 U3968 ( .A1(n4091), .A2(n7278), .ZN(n7279) );
  INV_X4 U3969 ( .A(n6728), .ZN(n6608) );
  NAND2_X2 U3970 ( .A1(net241770), .A2(net241771), .ZN(n4347) );
  NOR2_X2 U3971 ( .A1(net242655), .A2(net247632), .ZN(n3877) );
  NOR2_X4 U3972 ( .A1(n7400), .A2(n3878), .ZN(n7636) );
  INV_X4 U3973 ( .A(n3877), .ZN(n3878) );
  NOR2_X2 U3974 ( .A1(net242878), .A2(net247632), .ZN(n3879) );
  NOR2_X4 U3975 ( .A1(net242877), .A2(n3880), .ZN(n7393) );
  INV_X4 U3976 ( .A(n3879), .ZN(n3880) );
  NAND2_X2 U3977 ( .A1(b[9]), .A2(a[31]), .ZN(n3881) );
  NAND2_X2 U3978 ( .A1(n3882), .A2(n6935), .ZN(n7232) );
  INV_X4 U3979 ( .A(n3881), .ZN(n3882) );
  INV_X8 U3980 ( .A(b[7]), .ZN(net242655) );
  NAND2_X2 U3981 ( .A1(n7637), .A2(n7636), .ZN(n7638) );
  INV_X8 U3982 ( .A(b[8]), .ZN(net242878) );
  NAND2_X2 U3983 ( .A1(n7394), .A2(n7393), .ZN(n7395) );
  NAND2_X1 U3984 ( .A1(n4220), .A2(net242824), .ZN(n3885) );
  NAND2_X2 U3985 ( .A1(n3883), .A2(n3884), .ZN(n3886) );
  NAND2_X2 U3986 ( .A1(n3885), .A2(n3886), .ZN(n4218) );
  INV_X4 U3987 ( .A(n4220), .ZN(n3883) );
  INV_X1 U3988 ( .A(net242824), .ZN(n3884) );
  INV_X1 U3989 ( .A(n3888), .ZN(n3887) );
  OR2_X2 U3990 ( .A1(n4076), .A2(n7223), .ZN(n3908) );
  NAND2_X2 U3991 ( .A1(n6880), .A2(n6879), .ZN(net243275) );
  INV_X8 U3992 ( .A(n4045), .ZN(n4307) );
  OAI22_X4 U3993 ( .A1(net243996), .A2(net243997), .B1(net243998), .B2(
        net243785), .ZN(net243860) );
  NAND2_X2 U3994 ( .A1(n4328), .A2(net243582), .ZN(net243297) );
  INV_X4 U3995 ( .A(net243582), .ZN(net243635) );
  NAND2_X4 U3996 ( .A1(net243311), .A2(net243113), .ZN(net248040) );
  BUF_X4 U3997 ( .A(n6876), .Z(n4527) );
  INV_X1 U3998 ( .A(net247544), .ZN(net247545) );
  NAND2_X2 U3999 ( .A1(n5096), .A2(n5094), .ZN(n4999) );
  XNOR2_X2 U4000 ( .A(n8047), .B(n8046), .ZN(n4392) );
  NAND2_X1 U4001 ( .A1(n6148), .A2(n6147), .ZN(n6149) );
  INV_X4 U4002 ( .A(n4883), .ZN(n4496) );
  INV_X2 U4003 ( .A(net246273), .ZN(n4369) );
  NAND2_X1 U4004 ( .A1(n8328), .A2(n8327), .ZN(n8329) );
  INV_X2 U4005 ( .A(n7772), .ZN(n7775) );
  OAI21_X4 U4006 ( .B1(n5099), .B2(n5098), .A(n5097), .ZN(n5101) );
  INV_X8 U4007 ( .A(n6692), .ZN(n6725) );
  INV_X4 U4008 ( .A(net243723), .ZN(n3889) );
  INV_X8 U4009 ( .A(n3889), .ZN(n3890) );
  NAND2_X4 U4010 ( .A1(n6680), .A2(n6679), .ZN(n6682) );
  NAND2_X2 U4011 ( .A1(n6534), .A2(n6533), .ZN(n6680) );
  INV_X2 U4012 ( .A(n6156), .ZN(n6105) );
  NAND2_X2 U4013 ( .A1(net244063), .A2(net244062), .ZN(n3893) );
  NAND2_X4 U4014 ( .A1(n3891), .A2(n3892), .ZN(n3894) );
  NAND2_X4 U4015 ( .A1(n3893), .A2(n3894), .ZN(net244001) );
  INV_X8 U4016 ( .A(net244063), .ZN(n3891) );
  INV_X8 U4017 ( .A(net244062), .ZN(n3892) );
  INV_X8 U4018 ( .A(net243776), .ZN(net244063) );
  NAND2_X4 U4019 ( .A1(net244001), .A2(net243789), .ZN(net243784) );
  INV_X8 U4020 ( .A(net244001), .ZN(net247847) );
  INV_X8 U4021 ( .A(n6756), .ZN(n6960) );
  INV_X4 U4022 ( .A(net244063), .ZN(net248395) );
  NAND2_X4 U4023 ( .A1(net243775), .A2(net248395), .ZN(net243771) );
  AOI211_X1 U4024 ( .C1(n8107), .C2(net246974), .A(n8106), .B(n4267), .ZN(
        n8143) );
  NAND2_X4 U4025 ( .A1(net243185), .A2(net243186), .ZN(net243184) );
  NAND2_X2 U4026 ( .A1(n6030), .A2(n6033), .ZN(n6036) );
  NAND2_X1 U4027 ( .A1(net243268), .A2(n4353), .ZN(n7063) );
  XNOR2_X2 U4028 ( .A(n5044), .B(n5089), .ZN(n5121) );
  NAND2_X2 U4029 ( .A1(n5088), .A2(n5886), .ZN(n5044) );
  NOR2_X4 U4030 ( .A1(n5919), .A2(n5915), .ZN(n5916) );
  AOI21_X4 U4031 ( .B1(n5094), .B2(n5093), .A(n5095), .ZN(n5099) );
  NAND2_X4 U4032 ( .A1(n8346), .A2(n8345), .ZN(n8560) );
  XNOR2_X2 U4033 ( .A(n6079), .B(n6078), .ZN(n4457) );
  INV_X1 U4034 ( .A(n7478), .ZN(n4394) );
  XNOR2_X1 U4035 ( .A(n7567), .B(n3946), .ZN(n7711) );
  NOR2_X4 U4036 ( .A1(net242311), .A2(n4138), .ZN(net242376) );
  OAI21_X2 U4037 ( .B1(net248800), .B2(net245901), .A(net245902), .ZN(
        net245899) );
  BUF_X8 U4038 ( .A(n8772), .Z(n4426) );
  NAND2_X4 U4039 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  INV_X2 U4040 ( .A(out[3]), .ZN(n4151) );
  NAND2_X4 U4041 ( .A1(n8284), .A2(b[2]), .ZN(n8326) );
  OAI21_X2 U4042 ( .B1(n7474), .B2(n7473), .A(n7472), .ZN(n7475) );
  NOR2_X2 U4043 ( .A1(n7471), .A2(n7470), .ZN(n7474) );
  NOR2_X4 U4044 ( .A1(n4058), .A2(n4063), .ZN(n4062) );
  INV_X4 U4045 ( .A(n4068), .ZN(n4063) );
  INV_X4 U4046 ( .A(n3895), .ZN(n3896) );
  INV_X2 U4047 ( .A(n4525), .ZN(n7801) );
  OAI21_X2 U4048 ( .B1(n4525), .B2(n7806), .A(n7805), .ZN(n7807) );
  INV_X1 U4049 ( .A(n7298), .ZN(n3897) );
  INV_X4 U4050 ( .A(n7272), .ZN(n3898) );
  INV_X4 U4051 ( .A(n3898), .ZN(n3899) );
  OAI21_X4 U4052 ( .B1(net242607), .B2(net242606), .A(net242608), .ZN(n3903)
         );
  XNOR2_X2 U4053 ( .A(n3901), .B(n3900), .ZN(n7507) );
  INV_X32 U4054 ( .A(n7503), .ZN(n3900) );
  XNOR2_X2 U4055 ( .A(n7501), .B(n7500), .ZN(n3901) );
  NAND2_X2 U4056 ( .A1(n7696), .A2(n7697), .ZN(n7607) );
  OAI21_X2 U4057 ( .B1(n6805), .B2(n6806), .A(n6804), .ZN(n6808) );
  XNOR2_X2 U4058 ( .A(net241586), .B(net241063), .ZN(n3902) );
  OAI21_X2 U4059 ( .B1(net242607), .B2(net242606), .A(net242608), .ZN(
        net242605) );
  INV_X4 U4060 ( .A(net248357), .ZN(net245773) );
  OAI21_X2 U4061 ( .B1(net242604), .B2(net242603), .A(n3903), .ZN(net242303)
         );
  INV_X2 U4062 ( .A(n4396), .ZN(n5015) );
  XNOR2_X2 U4063 ( .A(n5139), .B(net248449), .ZN(n3904) );
  INV_X8 U4064 ( .A(n5002), .ZN(n5014) );
  INV_X2 U4065 ( .A(n8562), .ZN(n8754) );
  OAI21_X2 U4066 ( .B1(n8562), .B2(n8563), .A(n8561), .ZN(n8746) );
  XOR2_X1 U4067 ( .A(n7647), .B(n5643), .Z(n3905) );
  OAI21_X4 U4068 ( .B1(n4694), .B2(net246470), .A(n4693), .ZN(n4376) );
  INV_X8 U4069 ( .A(n4711), .ZN(n4713) );
  NOR2_X4 U4070 ( .A1(n5027), .A2(n5026), .ZN(n4911) );
  INV_X8 U4071 ( .A(n4928), .ZN(n4925) );
  OAI21_X4 U4072 ( .B1(n6340), .B2(n6339), .A(n6338), .ZN(n6466) );
  NAND2_X4 U4073 ( .A1(net245904), .A2(net245905), .ZN(net245893) );
  NAND2_X4 U4074 ( .A1(n6520), .A2(n6519), .ZN(n6325) );
  NAND2_X4 U4075 ( .A1(n5940), .A2(n5939), .ZN(n5083) );
  INV_X2 U4076 ( .A(net244665), .ZN(net247751) );
  AND2_X2 U4077 ( .A1(n6311), .A2(n6310), .ZN(n3906) );
  NAND2_X4 U4078 ( .A1(net244145), .A2(net244146), .ZN(net244143) );
  OAI21_X4 U4079 ( .B1(n4467), .B2(n6754), .A(n6753), .ZN(n6756) );
  INV_X4 U4080 ( .A(n6437), .ZN(n6674) );
  NAND2_X4 U4081 ( .A1(net243404), .A2(net243405), .ZN(n4341) );
  NAND2_X4 U4082 ( .A1(n6882), .A2(n6881), .ZN(net243404) );
  NAND2_X4 U4083 ( .A1(n6873), .A2(n6872), .ZN(net248780) );
  OAI21_X4 U4084 ( .B1(net243182), .B2(net243181), .A(net248703), .ZN(
        net248987) );
  AND2_X2 U4085 ( .A1(net242672), .A2(net242674), .ZN(n3907) );
  NAND2_X4 U4086 ( .A1(n7596), .A2(n7595), .ZN(n7288) );
  AND2_X2 U4087 ( .A1(net242811), .A2(net242813), .ZN(n3909) );
  INV_X1 U4088 ( .A(n7368), .ZN(n7577) );
  NAND2_X4 U4089 ( .A1(n8069), .A2(n8068), .ZN(n7702) );
  AND2_X2 U4090 ( .A1(n7862), .A2(n7861), .ZN(n3910) );
  XNOR2_X1 U4091 ( .A(n7641), .B(n7642), .ZN(n3911) );
  AND3_X4 U4092 ( .A1(n8085), .A2(n8084), .A3(n8083), .ZN(n3912) );
  INV_X4 U4093 ( .A(net240933), .ZN(n4271) );
  NAND2_X4 U4094 ( .A1(net240995), .A2(net240996), .ZN(net240994) );
  INV_X8 U4095 ( .A(net244284), .ZN(net247544) );
  BUF_X8 U4096 ( .A(net243995), .Z(net247563) );
  INV_X2 U4097 ( .A(n5057), .ZN(n4124) );
  NAND2_X1 U4098 ( .A1(net246541), .A2(net245422), .ZN(n3915) );
  NAND2_X4 U4099 ( .A1(n3913), .A2(n3914), .ZN(n3916) );
  NAND2_X2 U4100 ( .A1(n3915), .A2(n3916), .ZN(net247843) );
  INV_X4 U4101 ( .A(net246541), .ZN(n3913) );
  INV_X4 U4102 ( .A(net245422), .ZN(n3914) );
  NAND2_X2 U4103 ( .A1(net244066), .A2(net247563), .ZN(n3919) );
  NAND2_X4 U4104 ( .A1(n3917), .A2(n3918), .ZN(n3920) );
  NAND2_X4 U4105 ( .A1(n3919), .A2(n3920), .ZN(n4288) );
  INV_X4 U4106 ( .A(net244066), .ZN(n3917) );
  NAND2_X2 U4107 ( .A1(n4801), .A2(net248350), .ZN(n3923) );
  NAND2_X4 U4108 ( .A1(n3921), .A2(n3922), .ZN(n3924) );
  NAND2_X4 U4109 ( .A1(n3924), .A2(n3923), .ZN(net246250) );
  INV_X4 U4110 ( .A(n4801), .ZN(n3921) );
  INV_X4 U4111 ( .A(net248350), .ZN(n3922) );
  NAND2_X2 U4112 ( .A1(net245612), .A2(net244684), .ZN(n3927) );
  NAND2_X4 U4113 ( .A1(n3925), .A2(n3926), .ZN(n3928) );
  NAND2_X4 U4114 ( .A1(n3927), .A2(n3928), .ZN(net244562) );
  INV_X4 U4115 ( .A(net245612), .ZN(n3925) );
  INV_X1 U4116 ( .A(net244684), .ZN(n3926) );
  NAND2_X4 U4117 ( .A1(n3934), .A2(net246250), .ZN(n4874) );
  NAND2_X4 U4118 ( .A1(net246250), .A2(net246251), .ZN(net246117) );
  NAND2_X1 U4119 ( .A1(net246836), .A2(net246768), .ZN(net244684) );
  OAI21_X4 U4120 ( .B1(n7504), .B2(n7503), .A(n7502), .ZN(n7505) );
  NAND2_X2 U4121 ( .A1(n7501), .A2(n7500), .ZN(n7502) );
  NOR2_X2 U4122 ( .A1(n7501), .A2(n7500), .ZN(n7504) );
  BUF_X4 U4123 ( .A(n7996), .Z(n4423) );
  NAND2_X4 U4124 ( .A1(net241061), .A2(n8758), .ZN(net240996) );
  OAI21_X4 U4125 ( .B1(n7310), .B2(n7309), .A(n7308), .ZN(n7477) );
  INV_X4 U4126 ( .A(n4380), .ZN(n4381) );
  OAI21_X2 U4127 ( .B1(net241062), .B2(net241063), .A(net241064), .ZN(
        net241050) );
  NAND2_X4 U4128 ( .A1(b[31]), .A2(a[27]), .ZN(net246534) );
  INV_X4 U4129 ( .A(n7892), .ZN(n8145) );
  NOR2_X2 U4130 ( .A1(net241065), .A2(n8751), .ZN(net241062) );
  INV_X4 U4131 ( .A(net244144), .ZN(net244285) );
  NAND2_X4 U4132 ( .A1(net242320), .A2(net242321), .ZN(net242305) );
  NAND2_X4 U4133 ( .A1(n4567), .A2(net246778), .ZN(net245349) );
  NOR2_X4 U4134 ( .A1(n4060), .A2(n4062), .ZN(n4070) );
  AOI21_X4 U4135 ( .B1(n4268), .B2(net240929), .A(net240939), .ZN(net240937)
         );
  INV_X8 U4136 ( .A(net246433), .ZN(n4239) );
  NOR3_X4 U4137 ( .A1(n8107), .A2(net247632), .A3(n8281), .ZN(n8767) );
  NOR2_X2 U4138 ( .A1(net246836), .A2(n4572), .ZN(n5515) );
  NOR2_X2 U4139 ( .A1(net246878), .A2(net246782), .ZN(n5498) );
  NAND3_X2 U4140 ( .A1(n5568), .A2(n5567), .A3(n5566), .ZN(n5569) );
  INV_X16 U4141 ( .A(n5995), .ZN(n4544) );
  INV_X4 U4142 ( .A(b[27]), .ZN(net246876) );
  AOI21_X2 U4143 ( .B1(n4557), .B2(n6408), .A(n6123), .ZN(n6128) );
  NOR2_X1 U4144 ( .A1(n6122), .A2(n4533), .ZN(n6123) );
  INV_X1 U4145 ( .A(n7510), .ZN(n4460) );
  AOI21_X1 U4146 ( .B1(n4988), .B2(n4987), .A(n5107), .ZN(n4989) );
  OAI21_X2 U4147 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8441) );
  OAI21_X2 U4148 ( .B1(n8615), .B2(n8614), .A(n8613), .ZN(n8707) );
  OAI21_X2 U4149 ( .B1(n8619), .B2(n8618), .A(n8617), .ZN(n8705) );
  OAI21_X2 U4150 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8709) );
  OAI21_X2 U4151 ( .B1(n8501), .B2(n8500), .A(n8499), .ZN(n8503) );
  NOR2_X2 U4152 ( .A1(out[27]), .A2(n8810), .ZN(n8812) );
  NOR2_X2 U4153 ( .A1(n4428), .A2(n8729), .ZN(n8731) );
  AOI21_X1 U4154 ( .B1(n4428), .B2(n8729), .A(n8728), .ZN(n8732) );
  NOR2_X2 U4155 ( .A1(net246772), .A2(net246874), .ZN(n5500) );
  NOR3_X1 U4156 ( .A1(n5709), .A2(n5710), .A3(n5708), .ZN(n5655) );
  NOR2_X2 U4157 ( .A1(n5632), .A2(n5631), .ZN(n5657) );
  NOR2_X2 U4158 ( .A1(n5636), .A2(n5635), .ZN(n5656) );
  NOR2_X2 U4159 ( .A1(n5653), .A2(n5652), .ZN(n5654) );
  NOR2_X1 U4160 ( .A1(n5649), .A2(n5697), .ZN(n5650) );
  NOR2_X2 U4161 ( .A1(n5545), .A2(n5544), .ZN(n5608) );
  NOR3_X2 U4162 ( .A1(n5561), .A2(n5560), .A3(n5559), .ZN(n5607) );
  NOR2_X1 U4163 ( .A1(n6553), .A2(net247083), .ZN(n5177) );
  AOI21_X1 U4164 ( .B1(net246962), .B2(net246766), .A(n5187), .ZN(n5188) );
  NOR2_X1 U4165 ( .A1(n6901), .A2(net247083), .ZN(n5185) );
  NOR2_X1 U4166 ( .A1(n7029), .A2(net247083), .ZN(n5160) );
  NOR2_X2 U4167 ( .A1(n7240), .A2(net247083), .ZN(n5182) );
  NAND3_X2 U4168 ( .A1(n3982), .A2(n7421), .A3(n7420), .ZN(n8303) );
  INV_X4 U4169 ( .A(n7830), .ZN(n4532) );
  NAND2_X2 U4170 ( .A1(b[29]), .A2(net248517), .ZN(n7830) );
  NAND2_X2 U4171 ( .A1(n4496), .A2(net247817), .ZN(n4498) );
  NOR2_X2 U4172 ( .A1(n5422), .A2(n4572), .ZN(n4614) );
  INV_X4 U4173 ( .A(net240917), .ZN(net247059) );
  NOR2_X2 U4174 ( .A1(n6343), .A2(n6342), .ZN(n6345) );
  INV_X1 U4175 ( .A(n7530), .ZN(n4047) );
  INV_X4 U4176 ( .A(n4101), .ZN(n7927) );
  OAI21_X2 U4177 ( .B1(n7198), .B2(n7197), .A(n7196), .ZN(n7200) );
  NOR2_X1 U4178 ( .A1(n5107), .A2(n5872), .ZN(n5108) );
  AOI21_X2 U4179 ( .B1(n5106), .B2(n5105), .A(n5104), .ZN(n5109) );
  INV_X4 U4180 ( .A(n8358), .ZN(n4079) );
  INV_X4 U4181 ( .A(n7157), .ZN(n4077) );
  OAI21_X2 U4182 ( .B1(n7300), .B2(n7459), .A(n7457), .ZN(n7464) );
  INV_X4 U4183 ( .A(n8448), .ZN(n4374) );
  NOR2_X2 U4184 ( .A1(n6525), .A2(n6660), .ZN(n6663) );
  INV_X2 U4185 ( .A(n7597), .ZN(n4087) );
  OAI21_X2 U4186 ( .B1(n8603), .B2(n8602), .A(n8601), .ZN(n8713) );
  OAI21_X2 U4187 ( .B1(n8607), .B2(n8606), .A(n8605), .ZN(n8711) );
  OAI21_X2 U4188 ( .B1(n8599), .B2(n8598), .A(n8597), .ZN(n8715) );
  OAI21_X2 U4189 ( .B1(n7704), .B2(n4040), .A(n7703), .ZN(n8052) );
  OAI21_X2 U4190 ( .B1(n8583), .B2(n8582), .A(n8581), .ZN(n8736) );
  NOR2_X2 U4191 ( .A1(a[14]), .A2(net244239), .ZN(n5529) );
  NAND2_X1 U4192 ( .A1(net242610), .A2(net242609), .ZN(net242612) );
  NAND2_X2 U4193 ( .A1(net241040), .A2(net241018), .ZN(n8761) );
  NAND3_X2 U4194 ( .A1(net240812), .A2(net240813), .A3(net240761), .ZN(n4157)
         );
  NOR2_X1 U4195 ( .A1(net246766), .A2(net246868), .ZN(n5503) );
  NAND3_X1 U4196 ( .A1(n5696), .A2(n3905), .A3(n5695), .ZN(n5701) );
  NOR2_X2 U4197 ( .A1(n5694), .A2(n5693), .ZN(n5695) );
  NOR3_X2 U4198 ( .A1(n5698), .A2(n5770), .A3(n5697), .ZN(n5699) );
  NOR3_X2 U4199 ( .A1(n5605), .A2(n5604), .A3(n5769), .ZN(n5606) );
  NOR2_X1 U4200 ( .A1(n5770), .A2(n5765), .ZN(n5686) );
  NOR2_X1 U4201 ( .A1(n6398), .A2(net247083), .ZN(n5213) );
  NAND3_X2 U4202 ( .A1(n5340), .A2(a[31]), .A3(b[24]), .ZN(n4798) );
  AOI21_X2 U4203 ( .B1(n4561), .B2(n6280), .A(n6279), .ZN(n6285) );
  NOR2_X1 U4204 ( .A1(n6278), .A2(n8832), .ZN(n6279) );
  AOI21_X1 U4205 ( .B1(n8303), .B2(n4564), .A(n3995), .ZN(n7422) );
  NOR2_X1 U4206 ( .A1(n8833), .A2(n8832), .ZN(n8838) );
  AOI21_X2 U4207 ( .B1(n8792), .B2(n8791), .A(n4566), .ZN(n8793) );
  NOR2_X1 U4208 ( .A1(n1323), .A2(n8843), .ZN(n8844) );
  NOR2_X2 U4209 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  OAI21_X1 U4210 ( .B1(n5790), .B2(n4533), .A(n5789), .ZN(n5798) );
  AOI21_X2 U4211 ( .B1(n5242), .B2(n5241), .A(n4566), .ZN(n5243) );
  NOR2_X1 U4212 ( .A1(n5323), .A2(n4539), .ZN(n5324) );
  AOI21_X2 U4213 ( .B1(net245389), .B2(n5319), .A(n3996), .ZN(n5321) );
  INV_X8 U4214 ( .A(b[24]), .ZN(net246856) );
  AOI21_X2 U4215 ( .B1(n3977), .B2(n5480), .A(n5376), .ZN(n5377) );
  NOR2_X2 U4216 ( .A1(n5472), .A2(n4575), .ZN(n4620) );
  AOI21_X2 U4217 ( .B1(n4561), .B2(n5818), .A(n4655), .ZN(n4660) );
  NOR2_X1 U4218 ( .A1(n6122), .A2(n8832), .ZN(n4655) );
  NOR2_X1 U4219 ( .A1(n5993), .A2(n4537), .ZN(n6004) );
  NOR2_X2 U4220 ( .A1(n6117), .A2(n4580), .ZN(n6120) );
  OAI21_X1 U4221 ( .B1(n6272), .B2(n4531), .A(n6271), .ZN(n6289) );
  NOR2_X1 U4222 ( .A1(n6418), .A2(n4535), .ZN(n6288) );
  OAI21_X1 U4223 ( .B1(n6574), .B2(n4531), .A(n6573), .ZN(n6575) );
  NOR2_X1 U4224 ( .A1(n6705), .A2(n4537), .ZN(n6706) );
  NOR2_X2 U4225 ( .A1(n6713), .A2(n6712), .ZN(n6716) );
  AOI21_X1 U4226 ( .B1(n4555), .B2(n7256), .A(n3997), .ZN(n6914) );
  OAI21_X1 U4227 ( .B1(n6911), .B2(n4531), .A(n6910), .ZN(n6926) );
  NOR2_X1 U4228 ( .A1(n7255), .A2(n4535), .ZN(n7049) );
  NOR2_X1 U4229 ( .A1(n7047), .A2(n4531), .ZN(n7048) );
  NOR2_X1 U4230 ( .A1(n7418), .A2(n4535), .ZN(n7260) );
  OAI21_X1 U4231 ( .B1(n7255), .B2(n4531), .A(n7254), .ZN(n7261) );
  NOR2_X2 U4232 ( .A1(n7410), .A2(n7409), .ZN(n7413) );
  AOI21_X1 U4233 ( .B1(n4555), .B2(n8111), .A(n7656), .ZN(n7657) );
  OAI21_X1 U4234 ( .B1(n1386), .B2(n4566), .A(n7832), .ZN(n8109) );
  AOI21_X1 U4235 ( .B1(n4555), .B2(n8314), .A(n8112), .ZN(n7832) );
  NOR2_X2 U4236 ( .A1(n8290), .A2(n8289), .ZN(n8293) );
  OAI21_X1 U4237 ( .B1(n8313), .B2(n4531), .A(n8311), .ZN(n8317) );
  INV_X4 U4238 ( .A(n4545), .ZN(n4549) );
  INV_X4 U4239 ( .A(n8850), .ZN(n4540) );
  AOI21_X2 U4240 ( .B1(n5279), .B2(n5278), .A(n4547), .ZN(n5280) );
  NOR2_X2 U4241 ( .A1(net246874), .A2(net246970), .ZN(n5258) );
  OAI21_X2 U4242 ( .B1(b[27]), .B2(net247060), .A(n4550), .ZN(n5257) );
  NOR2_X2 U4243 ( .A1(net246832), .A2(net240784), .ZN(n5441) );
  OAI21_X2 U4244 ( .B1(b[20]), .B2(net247060), .A(n4550), .ZN(n5440) );
  NOR2_X2 U4245 ( .A1(n7490), .A2(n7491), .ZN(n7494) );
  NOR2_X2 U4246 ( .A1(n7507), .A2(n7508), .ZN(n7511) );
  NOR2_X2 U4247 ( .A1(n6626), .A2(n6625), .ZN(n6629) );
  NOR2_X2 U4248 ( .A1(n4433), .A2(n7517), .ZN(n7521) );
  NOR2_X2 U4249 ( .A1(n7538), .A2(n7537), .ZN(n7541) );
  NOR2_X2 U4250 ( .A1(n7486), .A2(n7485), .ZN(n7488) );
  OAI21_X2 U4251 ( .B1(n7548), .B2(n7547), .A(n3976), .ZN(n7549) );
  INV_X4 U4252 ( .A(n7959), .ZN(n4049) );
  INV_X2 U4253 ( .A(n7137), .ZN(n4389) );
  INV_X4 U4254 ( .A(n6481), .ZN(n6479) );
  NAND2_X2 U4255 ( .A1(n6488), .A2(n6487), .ZN(n6490) );
  AOI21_X2 U4256 ( .B1(n5873), .B2(n5872), .A(n5871), .ZN(n5875) );
  NOR2_X2 U4257 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  AOI21_X2 U4258 ( .B1(n6495), .B2(n6494), .A(n6497), .ZN(n6501) );
  OAI21_X2 U4259 ( .B1(n8000), .B2(n7999), .A(n7998), .ZN(n8002) );
  NOR2_X2 U4260 ( .A1(n4423), .A2(n7997), .ZN(n8000) );
  INV_X4 U4261 ( .A(n7997), .ZN(n4088) );
  INV_X4 U4262 ( .A(n8398), .ZN(n4055) );
  NAND2_X2 U4263 ( .A1(n6329), .A2(n6328), .ZN(n6326) );
  INV_X4 U4264 ( .A(n7167), .ZN(n4424) );
  OAI21_X2 U4265 ( .B1(n7455), .B2(n7454), .A(n7453), .ZN(n7456) );
  NOR2_X2 U4266 ( .A1(n8386), .A2(n8385), .ZN(n8389) );
  OAI21_X2 U4267 ( .B1(n8627), .B2(n8626), .A(n8625), .ZN(n8701) );
  OAI21_X2 U4268 ( .B1(n8631), .B2(n8630), .A(n8629), .ZN(n8699) );
  OAI21_X2 U4269 ( .B1(n8623), .B2(n8622), .A(n8621), .ZN(n8703) );
  INV_X4 U4270 ( .A(n6220), .ZN(n6224) );
  OAI21_X2 U4271 ( .B1(n6162), .B2(n6161), .A(n6160), .ZN(net244374) );
  NOR3_X2 U4272 ( .A1(n6162), .A2(n6160), .A3(n6161), .ZN(net244373) );
  NAND2_X2 U4273 ( .A1(n7090), .A2(n7091), .ZN(n7094) );
  NAND2_X2 U4274 ( .A1(net244077), .A2(net244075), .ZN(net244073) );
  NAND2_X2 U4275 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  OAI21_X2 U4276 ( .B1(n4816), .B2(n4814), .A(n4813), .ZN(n4818) );
  NAND3_X2 U4277 ( .A1(n6737), .A2(n6736), .A3(n6738), .ZN(n6675) );
  OAI21_X2 U4278 ( .B1(n8591), .B2(n8590), .A(n8589), .ZN(n8719) );
  OAI21_X2 U4279 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8717) );
  AOI21_X2 U4280 ( .B1(n8587), .B2(n8586), .A(n8585), .ZN(n8721) );
  INV_X4 U4281 ( .A(net246886), .ZN(net246882) );
  NOR2_X2 U4282 ( .A1(net243770), .A2(n4183), .ZN(net243774) );
  INV_X4 U4283 ( .A(n6601), .ZN(n6865) );
  NOR2_X2 U4284 ( .A1(n8058), .A2(n8057), .ZN(n8061) );
  NOR2_X2 U4285 ( .A1(n8536), .A2(n8535), .ZN(n8528) );
  OAI21_X2 U4286 ( .B1(n4286), .B2(n4073), .A(net244674), .ZN(n4285) );
  INV_X4 U4287 ( .A(n3890), .ZN(n4186) );
  NAND2_X2 U4288 ( .A1(net243106), .A2(net243119), .ZN(n4343) );
  NAND2_X2 U4289 ( .A1(n8494), .A2(n8173), .ZN(n8046) );
  NOR2_X2 U4290 ( .A1(n3929), .A2(n4180), .ZN(net246488) );
  AOI21_X2 U4291 ( .B1(n6246), .B2(n6310), .A(n6312), .ZN(n6251) );
  INV_X4 U4292 ( .A(net248371), .ZN(net243757) );
  NAND2_X2 U4293 ( .A1(n6936), .A2(net243288), .ZN(net243286) );
  OAI21_X2 U4294 ( .B1(n8575), .B2(n8574), .A(n8573), .ZN(n8740) );
  NAND3_X2 U4295 ( .A1(n5546), .A2(n5623), .A3(n5621), .ZN(n5539) );
  NAND3_X2 U4296 ( .A1(n5551), .A2(n5614), .A3(n5616), .ZN(n5555) );
  NOR2_X2 U4297 ( .A1(a[16]), .A2(net244627), .ZN(n5525) );
  OAI21_X2 U4298 ( .B1(a[30]), .B2(net246790), .A(net248516), .ZN(net246530)
         );
  INV_X4 U4299 ( .A(net246467), .ZN(net247795) );
  INV_X4 U4300 ( .A(net245955), .ZN(net246081) );
  OAI21_X2 U4301 ( .B1(n8559), .B2(n8558), .A(n8557), .ZN(n8748) );
  NOR2_X2 U4302 ( .A1(n5694), .A2(n5692), .ZN(n5647) );
  NAND3_X2 U4303 ( .A1(n5579), .A2(n5578), .A3(n5577), .ZN(n5649) );
  NOR2_X2 U4304 ( .A1(net246788), .A2(n4569), .ZN(n5496) );
  NAND2_X1 U4305 ( .A1(b[23]), .A2(net246786), .ZN(n4876) );
  NAND2_X2 U4306 ( .A1(net243362), .A2(net243361), .ZN(n4179) );
  INV_X4 U4307 ( .A(n7227), .ZN(n4090) );
  OAI21_X2 U4308 ( .B1(net242672), .B2(net242673), .A(net242674), .ZN(
        net242669) );
  INV_X4 U4309 ( .A(net241831), .ZN(net242066) );
  NOR2_X1 U4310 ( .A1(n8289), .A2(n8298), .ZN(n5169) );
  NOR2_X1 U4311 ( .A1(n8773), .A2(n8298), .ZN(n5187) );
  NOR2_X2 U4312 ( .A1(n5945), .A2(n5946), .ZN(n4053) );
  INV_X4 U4313 ( .A(net243645), .ZN(net243639) );
  NOR2_X1 U4314 ( .A1(net246812), .A2(net247083), .ZN(n5987) );
  NAND3_X2 U4315 ( .A1(n6283), .A2(n6282), .A3(n6281), .ZN(n7247) );
  INV_X4 U4316 ( .A(n8258), .ZN(n8259) );
  INV_X8 U4317 ( .A(n8796), .ZN(n4560) );
  NAND3_X1 U4318 ( .A1(n6919), .A2(n6918), .A3(n6917), .ZN(n8118) );
  NOR2_X2 U4319 ( .A1(net246956), .A2(n8773), .ZN(n8300) );
  NOR2_X1 U4320 ( .A1(n4576), .A2(net247083), .ZN(n8296) );
  NAND2_X2 U4321 ( .A1(n8765), .A2(n8764), .ZN(net240975) );
  NOR2_X2 U4322 ( .A1(net240982), .A2(net240956), .ZN(net240981) );
  NOR3_X2 U4323 ( .A1(n5771), .A2(n5770), .A3(n5769), .ZN(n5772) );
  NOR2_X1 U4324 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  INV_X16 U4325 ( .A(a[25]), .ZN(net246764) );
  INV_X4 U4326 ( .A(net248925), .ZN(net246260) );
  NOR2_X1 U4327 ( .A1(net240839), .A2(net247083), .ZN(n4629) );
  INV_X8 U4328 ( .A(a[21]), .ZN(n4573) );
  NAND3_X2 U4329 ( .A1(n5997), .A2(n7038), .A3(n5996), .ZN(n6913) );
  INV_X4 U4330 ( .A(net243376), .ZN(net243373) );
  NOR2_X1 U4331 ( .A1(net246804), .A2(net247083), .ZN(n6124) );
  NAND3_X2 U4332 ( .A1(n6411), .A2(n6410), .A3(n6409), .ZN(n7419) );
  OAI21_X2 U4333 ( .B1(net246956), .B2(n7842), .A(n7044), .ZN(n7415) );
  NOR2_X1 U4334 ( .A1(n8786), .A2(n4569), .ZN(n8112) );
  NOR2_X1 U4335 ( .A1(net246812), .A2(n4357), .ZN(n4358) );
  AOI21_X2 U4336 ( .B1(n5716), .B2(n5715), .A(ALUCtrl[2]), .ZN(n5719) );
  NOR2_X2 U4337 ( .A1(n5671), .A2(n5670), .ZN(n5689) );
  NOR2_X2 U4338 ( .A1(n5693), .A2(n5687), .ZN(n5688) );
  NOR2_X2 U4339 ( .A1(n5661), .A2(n5660), .ZN(n5690) );
  NOR2_X1 U4340 ( .A1(n5780), .A2(net244867), .ZN(n5781) );
  NOR2_X2 U4341 ( .A1(n5779), .A2(n5778), .ZN(n5782) );
  OAI21_X1 U4342 ( .B1(n5270), .B2(net245318), .A(n5269), .ZN(n5301) );
  NOR2_X2 U4343 ( .A1(b[26]), .A2(net246766), .ZN(n5287) );
  INV_X16 U4344 ( .A(n3987), .ZN(n4545) );
  NOR2_X1 U4345 ( .A1(net246924), .A2(net244841), .ZN(n4670) );
  NOR2_X2 U4346 ( .A1(n5365), .A2(net246750), .ZN(n4608) );
  NOR2_X2 U4347 ( .A1(n5845), .A2(n4577), .ZN(n4626) );
  NOR2_X2 U4348 ( .A1(n6399), .A2(n6398), .ZN(n6402) );
  NOR2_X2 U4349 ( .A1(n7030), .A2(n7029), .ZN(n7033) );
  NOR2_X2 U4350 ( .A1(n7843), .A2(n7842), .ZN(n7846) );
  OAI21_X1 U4351 ( .B1(n1323), .B2(n4566), .A(n8786), .ZN(n8787) );
  NOR2_X2 U4352 ( .A1(n8845), .A2(n8844), .ZN(n8846) );
  NOR2_X1 U4353 ( .A1(n8851), .A2(n4541), .ZN(n8852) );
  AOI21_X2 U4354 ( .B1(n8827), .B2(net240852), .A(n8826), .ZN(n8829) );
  NOR2_X2 U4355 ( .A1(n8827), .A2(net240852), .ZN(n8828) );
  OAI21_X1 U4356 ( .B1(n5800), .B2(n4535), .A(n5799), .ZN(n5802) );
  OAI21_X2 U4357 ( .B1(n5798), .B2(n5797), .A(n8842), .ZN(n5799) );
  OAI21_X1 U4358 ( .B1(n5796), .B2(n8115), .A(n5795), .ZN(n5797) );
  AOI21_X1 U4359 ( .B1(net240784), .B2(net247048), .A(net246918), .ZN(n5801)
         );
  NOR2_X2 U4360 ( .A1(n5808), .A2(n4541), .ZN(n5809) );
  NOR3_X1 U4361 ( .A1(net245388), .A2(n3978), .A3(net247060), .ZN(n5251) );
  NAND3_X1 U4362 ( .A1(n4264), .A2(net245388), .A3(n3978), .ZN(net245474) );
  NOR2_X2 U4363 ( .A1(n4541), .A2(n5748), .ZN(n5238) );
  NOR2_X1 U4364 ( .A1(net247044), .A2(n5236), .ZN(n5237) );
  NOR2_X1 U4365 ( .A1(n4569), .A2(net246970), .ZN(net245524) );
  OAI21_X2 U4366 ( .B1(b[29]), .B2(net247060), .A(n4550), .ZN(net245525) );
  NOR2_X2 U4367 ( .A1(n4541), .A2(n5678), .ZN(n5209) );
  INV_X16 U4368 ( .A(net247044), .ZN(net240782) );
  NOR2_X1 U4369 ( .A1(net246878), .A2(net247060), .ZN(n5196) );
  NOR2_X1 U4370 ( .A1(net245541), .A2(net247044), .ZN(n5199) );
  NOR2_X2 U4371 ( .A1(net246868), .A2(net246970), .ZN(n5286) );
  OAI21_X2 U4372 ( .B1(b[26]), .B2(net247060), .A(n4550), .ZN(n5285) );
  NOR2_X2 U4373 ( .A1(b[25]), .A2(net247060), .ZN(n5330) );
  NOR2_X1 U4374 ( .A1(n5322), .A2(n4537), .ZN(n5325) );
  NOR2_X1 U4375 ( .A1(net245369), .A2(net247044), .ZN(n5334) );
  NOR2_X2 U4376 ( .A1(net246970), .A2(net246856), .ZN(net245359) );
  OAI21_X2 U4377 ( .B1(b[24]), .B2(net247060), .A(n4550), .ZN(n5341) );
  NOR2_X2 U4378 ( .A1(b[23]), .A2(net247060), .ZN(n5369) );
  NOR2_X1 U4379 ( .A1(n4541), .A2(n5672), .ZN(n5367) );
  NOR2_X1 U4380 ( .A1(n5385), .A2(net247048), .ZN(n5386) );
  NOR2_X1 U4381 ( .A1(n6037), .A2(net247044), .ZN(n5387) );
  NOR2_X2 U4382 ( .A1(b[22]), .A2(net247060), .ZN(n5410) );
  AOI21_X2 U4383 ( .B1(n5407), .B2(n5406), .A(n4547), .ZN(n5408) );
  NOR2_X1 U4384 ( .A1(n6322), .A2(net247044), .ZN(n5413) );
  NOR2_X2 U4385 ( .A1(net246838), .A2(net240784), .ZN(net245266) );
  OAI21_X1 U4386 ( .B1(net246836), .B2(net247060), .A(n4550), .ZN(n5418) );
  NOR2_X2 U4387 ( .A1(n4145), .A2(net240784), .ZN(net245207) );
  OAI21_X2 U4388 ( .B1(b[19]), .B2(net247060), .A(n4550), .ZN(n5466) );
  NOR2_X2 U4389 ( .A1(b[18]), .A2(net247060), .ZN(n5833) );
  NOR2_X1 U4390 ( .A1(n7767), .A2(net247044), .ZN(n5838) );
  NOR2_X2 U4391 ( .A1(b[17]), .A2(net247060), .ZN(n5854) );
  NOR2_X1 U4392 ( .A1(n8182), .A2(net247044), .ZN(n5858) );
  NOR2_X2 U4393 ( .A1(b[16]), .A2(net247060), .ZN(n4675) );
  AOI21_X1 U4394 ( .B1(n4672), .B2(n4671), .A(n4547), .ZN(n4673) );
  NOR2_X1 U4395 ( .A1(n8729), .A2(net247044), .ZN(n5151) );
  OAI21_X1 U4396 ( .B1(n6007), .B2(n4546), .A(n6006), .ZN(n6008) );
  NOR2_X1 U4397 ( .A1(n6002), .A2(n4535), .ZN(n6003) );
  OAI21_X1 U4398 ( .B1(n6139), .B2(n4546), .A(n6138), .ZN(n6140) );
  OAI21_X1 U4399 ( .B1(n6291), .B2(n4546), .A(n6290), .ZN(n6292) );
  NOR2_X1 U4400 ( .A1(n6286), .A2(n4537), .ZN(n6287) );
  OAI21_X1 U4401 ( .B1(n6421), .B2(n4546), .A(n6420), .ZN(n6422) );
  OAI21_X1 U4402 ( .B1(n6578), .B2(n4546), .A(n6577), .ZN(n6579) );
  OAI21_X1 U4403 ( .B1(n6571), .B2(n4535), .A(n6570), .ZN(n6576) );
  AOI21_X1 U4404 ( .B1(n6708), .B2(n6707), .A(n4547), .ZN(n6709) );
  AOI21_X1 U4405 ( .B1(n8842), .B2(n6696), .A(n6695), .ZN(n6708) );
  NOR2_X1 U4406 ( .A1(n6694), .A2(n4539), .ZN(n6695) );
  NOR2_X1 U4407 ( .A1(n6901), .A2(net247044), .ZN(n6690) );
  OAI21_X1 U4408 ( .B1(n6901), .B2(net247048), .A(n6719), .ZN(n6720) );
  OAI21_X1 U4409 ( .B1(n6928), .B2(n4546), .A(n6927), .ZN(n6929) );
  OAI21_X1 U4410 ( .B1(n7047), .B2(n4535), .A(n6924), .ZN(n6925) );
  OAI21_X1 U4411 ( .B1(n7052), .B2(n4546), .A(n7051), .ZN(n7053) );
  OAI21_X1 U4412 ( .B1(n7263), .B2(n4546), .A(n7262), .ZN(n7264) );
  NOR3_X2 U4413 ( .A1(n7261), .A2(n7260), .A3(n7259), .ZN(n7263) );
  NOR2_X1 U4414 ( .A1(n3984), .A2(n4539), .ZN(n7259) );
  OAI21_X1 U4415 ( .B1(n7429), .B2(n4546), .A(n7428), .ZN(n7430) );
  OAI21_X1 U4416 ( .B1(n7672), .B2(n4546), .A(n7671), .ZN(n7673) );
  NOR2_X2 U4417 ( .A1(n7670), .A2(n7669), .ZN(n7672) );
  OAI21_X1 U4418 ( .B1(n7667), .B2(n4535), .A(n7666), .ZN(n7670) );
  AOI21_X1 U4419 ( .B1(n7838), .B2(n7837), .A(n4547), .ZN(n7839) );
  NOR2_X1 U4420 ( .A1(n7834), .A2(n4539), .ZN(n7835) );
  NOR2_X1 U4421 ( .A1(n8130), .A2(net247044), .ZN(n7822) );
  OAI21_X1 U4422 ( .B1(n8130), .B2(net247049), .A(n7849), .ZN(n7850) );
  INV_X4 U4423 ( .A(n8280), .ZN(n8107) );
  NOR2_X1 U4424 ( .A1(n8289), .A2(net247044), .ZN(n8106) );
  AOI21_X1 U4425 ( .B1(n8127), .B2(n8126), .A(n4547), .ZN(n8128) );
  AOI21_X1 U4426 ( .B1(n8125), .B2(n8309), .A(n8124), .ZN(n8126) );
  NOR2_X1 U4427 ( .A1(n8123), .A2(n4537), .ZN(n8124) );
  OAI21_X1 U4428 ( .B1(n8289), .B2(net247049), .A(n8138), .ZN(n8139) );
  OAI21_X1 U4429 ( .B1(n8320), .B2(n4546), .A(n8319), .ZN(n8321) );
  NOR2_X1 U4430 ( .A1(n8315), .A2(n4535), .ZN(n8316) );
  OAI21_X1 U4431 ( .B1(b[0]), .B2(net247060), .A(n4550), .ZN(net240915) );
  AOI21_X1 U4432 ( .B1(n4261), .B2(net246970), .A(n4262), .ZN(n4260) );
  NOR2_X2 U4433 ( .A1(n5263), .A2(n5262), .ZN(n5283) );
  AOI21_X2 U4434 ( .B1(n4552), .B2(n5463), .A(n5462), .ZN(n5464) );
  AOI21_X2 U4435 ( .B1(n5461), .B2(n5460), .A(n4547), .ZN(n5462) );
  NOR2_X2 U4436 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  NOR2_X2 U4437 ( .A1(n8862), .A2(net240772), .ZN(n8868) );
  INV_X16 U4438 ( .A(n4533), .ZN(n4562) );
  INV_X8 U4439 ( .A(a[28]), .ZN(net246782) );
  INV_X4 U4440 ( .A(net246782), .ZN(net246778) );
  INV_X16 U4441 ( .A(a[22]), .ZN(n4571) );
  INV_X8 U4442 ( .A(n4550), .ZN(n4551) );
  INV_X16 U4443 ( .A(a[20]), .ZN(n4574) );
  AND2_X4 U4444 ( .A1(b[27]), .A2(a[30]), .ZN(n3929) );
  AND2_X4 U4445 ( .A1(b[26]), .A2(net246772), .ZN(n3930) );
  INV_X16 U4446 ( .A(b[25]), .ZN(net246862) );
  AND2_X4 U4447 ( .A1(net240913), .A2(net246812), .ZN(n3931) );
  INV_X16 U4448 ( .A(n716), .ZN(n4563) );
  AND2_X2 U4449 ( .A1(n4765), .A2(n4764), .ZN(n3932) );
  INV_X4 U4450 ( .A(n4036), .ZN(net249274) );
  AND2_X4 U4451 ( .A1(a[23]), .A2(b[27]), .ZN(n3933) );
  AND2_X4 U4452 ( .A1(b[25]), .A2(a[28]), .ZN(n3934) );
  INV_X16 U4453 ( .A(b[22]), .ZN(net246844) );
  AND2_X2 U4454 ( .A1(a[19]), .A2(b[26]), .ZN(n3935) );
  AND2_X2 U4455 ( .A1(n6445), .A2(n6444), .ZN(n3936) );
  OR2_X2 U4456 ( .A1(out[6]), .A2(n3959), .ZN(n3937) );
  OR2_X2 U4457 ( .A1(out[8]), .A2(n3960), .ZN(n3938) );
  INV_X4 U4458 ( .A(b[17]), .ZN(n4570) );
  AND2_X4 U4459 ( .A1(a[21]), .A2(b[22]), .ZN(n3939) );
  AND2_X2 U4460 ( .A1(n7720), .A2(n7719), .ZN(n3940) );
  AND2_X2 U4461 ( .A1(n8196), .A2(n8195), .ZN(n3941) );
  OR2_X2 U4462 ( .A1(out[13]), .A2(n3972), .ZN(n3942) );
  INV_X16 U4463 ( .A(n5990), .ZN(n4556) );
  INV_X16 U4464 ( .A(n4556), .ZN(n4555) );
  INV_X16 U4465 ( .A(n4536), .ZN(n4537) );
  INV_X4 U4466 ( .A(n8848), .ZN(n4536) );
  OR2_X2 U4467 ( .A1(n7870), .A2(n7869), .ZN(n3943) );
  INV_X16 U4468 ( .A(b[29]), .ZN(n4568) );
  OR2_X2 U4469 ( .A1(net241070), .A2(net241071), .ZN(n3944) );
  OR2_X1 U4470 ( .A1(n7274), .A2(n7223), .ZN(n3945) );
  INV_X4 U4471 ( .A(net245963), .ZN(net249300) );
  XOR2_X2 U4472 ( .A(n7566), .B(n7763), .Z(n3946) );
  AND2_X2 U4473 ( .A1(n8554), .A2(n8553), .ZN(n3947) );
  INV_X4 U4474 ( .A(n7184), .ZN(n4108) );
  AND3_X4 U4475 ( .A1(n8182), .A2(n8181), .A3(n8180), .ZN(n3948) );
  AND3_X4 U4476 ( .A1(n7442), .A2(net242594), .A3(net242595), .ZN(n3949) );
  AND2_X4 U4477 ( .A1(n5955), .A2(n5954), .ZN(n3950) );
  OR3_X2 U4478 ( .A1(net242580), .A2(net242581), .A3(n7450), .ZN(n3951) );
  OR2_X2 U4479 ( .A1(out[2]), .A2(n4149), .ZN(n3952) );
  OR2_X2 U4480 ( .A1(n4903), .A2(n4859), .ZN(n3953) );
  AND2_X2 U4481 ( .A1(n4876), .A2(n4875), .ZN(n3954) );
  OR2_X2 U4482 ( .A1(n4815), .A2(n4767), .ZN(n3955) );
  AND2_X4 U4483 ( .A1(a[21]), .A2(b[29]), .ZN(n3956) );
  AND2_X4 U4484 ( .A1(b[22]), .A2(net246786), .ZN(n3957) );
  AND2_X2 U4485 ( .A1(a[10]), .A2(net248516), .ZN(n3958) );
  OR2_X2 U4486 ( .A1(out[7]), .A2(n3938), .ZN(n3959) );
  OR2_X2 U4487 ( .A1(out[9]), .A2(n4152), .ZN(n3960) );
  OR2_X4 U4488 ( .A1(n6446), .A2(n6624), .ZN(n3961) );
  INV_X4 U4489 ( .A(n5908), .ZN(n4488) );
  OR2_X1 U4490 ( .A1(n6341), .A2(n6174), .ZN(n3962) );
  OR2_X1 U4491 ( .A1(n7484), .A2(n7318), .ZN(n3963) );
  INV_X2 U4492 ( .A(net246111), .ZN(net246108) );
  OR2_X2 U4493 ( .A1(out[5]), .A2(n3937), .ZN(n3964) );
  AND2_X4 U4494 ( .A1(b[19]), .A2(net246772), .ZN(n3965) );
  AND2_X4 U4495 ( .A1(b[21]), .A2(a[30]), .ZN(n3966) );
  AND2_X4 U4496 ( .A1(b[18]), .A2(net246766), .ZN(n3967) );
  AND2_X4 U4497 ( .A1(a[16]), .A2(b[27]), .ZN(n3968) );
  INV_X4 U4498 ( .A(net245962), .ZN(net248207) );
  AND2_X2 U4499 ( .A1(a[18]), .A2(b[25]), .ZN(n3969) );
  AND2_X2 U4500 ( .A1(a[8]), .A2(net246880), .ZN(n3970) );
  OR2_X2 U4501 ( .A1(out[12]), .A2(n3942), .ZN(n3971) );
  OR2_X2 U4502 ( .A1(out[14]), .A2(n4155), .ZN(n3972) );
  INV_X4 U4503 ( .A(net244704), .ZN(net247168) );
  OR2_X4 U4504 ( .A1(n7721), .A2(n7909), .ZN(n3973) );
  OR2_X4 U4505 ( .A1(n8197), .A2(n8348), .ZN(n3974) );
  INV_X4 U4506 ( .A(net244273), .ZN(net248029) );
  AND2_X4 U4507 ( .A1(a[2]), .A2(net246904), .ZN(n3975) );
  INV_X4 U4508 ( .A(n7274), .ZN(n4091) );
  AND2_X2 U4509 ( .A1(a[14]), .A2(b[23]), .ZN(n3976) );
  AND2_X4 U4510 ( .A1(net246908), .A2(n4569), .ZN(n3977) );
  INV_X16 U4511 ( .A(net247082), .ZN(net247083) );
  INV_X16 U4512 ( .A(net241542), .ZN(net247082) );
  AND2_X4 U4513 ( .A1(net246916), .A2(a[30]), .ZN(n3978) );
  AND2_X4 U4514 ( .A1(a[18]), .A2(b[16]), .ZN(n3979) );
  INV_X2 U4515 ( .A(net245318), .ZN(net245389) );
  AND2_X4 U4516 ( .A1(net246760), .A2(b[10]), .ZN(n3980) );
  AND2_X2 U4517 ( .A1(b[9]), .A2(net246754), .ZN(n3981) );
  OR2_X4 U4518 ( .A1(net246956), .A2(n7648), .ZN(n3982) );
  AND2_X2 U4519 ( .A1(b[13]), .A2(net246754), .ZN(n3983) );
  INV_X4 U4520 ( .A(n4560), .ZN(n4559) );
  AND3_X4 U4521 ( .A1(n7042), .A2(n7041), .A3(n7040), .ZN(n3984) );
  AND3_X4 U4522 ( .A1(n5704), .A2(n5703), .A3(n5702), .ZN(n3985) );
  AND2_X4 U4523 ( .A1(n7423), .A2(n7422), .ZN(n3986) );
  NAND2_X1 U4524 ( .A1(b[6]), .A2(net246772), .ZN(net241039) );
  AND2_X4 U4525 ( .A1(n4670), .A2(n4669), .ZN(n3987) );
  OR2_X2 U4526 ( .A1(net246878), .A2(a[28]), .ZN(n3988) );
  OR2_X2 U4527 ( .A1(a[22]), .A2(b[22]), .ZN(n3989) );
  OR2_X4 U4528 ( .A1(a[18]), .A2(b[18]), .ZN(n3990) );
  OR2_X2 U4529 ( .A1(a[16]), .A2(b[16]), .ZN(n3991) );
  INV_X8 U4530 ( .A(n8781), .ZN(n4553) );
  INV_X16 U4531 ( .A(n4553), .ZN(n4552) );
  AND2_X2 U4532 ( .A1(n6697), .A2(n4565), .ZN(n3992) );
  OR2_X4 U4533 ( .A1(net246836), .A2(a[21]), .ZN(n3993) );
  AND2_X4 U4534 ( .A1(b[2]), .A2(a[31]), .ZN(n3994) );
  AND2_X2 U4535 ( .A1(n4555), .A2(n8305), .ZN(n3995) );
  AND3_X2 U4536 ( .A1(net246962), .A2(net245393), .A3(net246908), .ZN(n3996)
         );
  AND2_X2 U4537 ( .A1(n6913), .A2(n4565), .ZN(n3997) );
  AND2_X2 U4538 ( .A1(n8837), .A2(n4565), .ZN(n3998) );
  INV_X16 U4539 ( .A(n890), .ZN(net246966) );
  OR2_X4 U4540 ( .A1(net244627), .A2(net240784), .ZN(n3999) );
  INV_X16 U4541 ( .A(n4534), .ZN(n4535) );
  INV_X4 U4542 ( .A(n8806), .ZN(n4534) );
  INV_X16 U4543 ( .A(n4530), .ZN(n4531) );
  INV_X4 U4544 ( .A(n8312), .ZN(n4530) );
  OR2_X4 U4545 ( .A1(net246862), .A2(net240784), .ZN(n4000) );
  OR2_X4 U4546 ( .A1(net246844), .A2(net240784), .ZN(n4001) );
  OR2_X4 U4547 ( .A1(n4570), .A2(net240784), .ZN(n4002) );
  OR2_X4 U4548 ( .A1(n4323), .A2(net246970), .ZN(n4003) );
  INV_X1 U4549 ( .A(n4533), .ZN(n6564) );
  OR2_X2 U4550 ( .A1(net246850), .A2(net240784), .ZN(n4004) );
  OR2_X4 U4551 ( .A1(net244808), .A2(net240784), .ZN(n4005) );
  INV_X16 U4552 ( .A(n4538), .ZN(n4539) );
  INV_X4 U4553 ( .A(n8804), .ZN(n4538) );
  INV_X16 U4554 ( .A(net240784), .ZN(net246974) );
  INV_X2 U4555 ( .A(n4219), .ZN(n4006) );
  OAI211_X2 U4556 ( .C1(n3911), .C2(net246970), .A(net247049), .B(n7643), .ZN(
        n7644) );
  AOI21_X2 U4557 ( .B1(n6710), .B2(n6725), .A(n6709), .ZN(n6723) );
  NAND2_X2 U4558 ( .A1(n7229), .A2(n7230), .ZN(net242674) );
  NAND2_X2 U4559 ( .A1(net243765), .A2(n4289), .ZN(net243754) );
  XNOR2_X2 U4560 ( .A(net244270), .B(net248551), .ZN(n4007) );
  NAND2_X1 U4561 ( .A1(n4497), .A2(n4498), .ZN(n4008) );
  CLKBUF_X2 U4562 ( .A(net243765), .Z(n4009) );
  NOR2_X2 U4563 ( .A1(out[4]), .A2(n3964), .ZN(n4150) );
  OAI211_X2 U4564 ( .C1(n4426), .C2(net246970), .A(net247048), .B(n8283), .ZN(
        n8284) );
  NAND2_X4 U4565 ( .A1(n7707), .A2(n7706), .ZN(n7593) );
  NOR2_X2 U4566 ( .A1(n8426), .A2(n8425), .ZN(n8429) );
  NAND2_X1 U4567 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  NOR2_X1 U4568 ( .A1(n8435), .A2(n8436), .ZN(n8439) );
  NAND2_X1 U4569 ( .A1(n8436), .A2(n8435), .ZN(n8437) );
  XNOR2_X2 U4570 ( .A(n5928), .B(n5927), .ZN(n4010) );
  NOR2_X4 U4571 ( .A1(n6682), .A2(n6681), .ZN(n4075) );
  INV_X8 U4572 ( .A(net242602), .ZN(net242597) );
  NAND2_X2 U4573 ( .A1(n7620), .A2(net242402), .ZN(n7621) );
  NAND2_X4 U4574 ( .A1(n4099), .A2(n3899), .ZN(n7620) );
  INV_X1 U4575 ( .A(n7175), .ZN(n4011) );
  INV_X2 U4576 ( .A(n4011), .ZN(n4012) );
  XNOR2_X2 U4577 ( .A(n7002), .B(n7174), .ZN(n4013) );
  XNOR2_X2 U4578 ( .A(n6659), .B(n6823), .ZN(n4014) );
  NAND2_X4 U4579 ( .A1(n4483), .A2(n4482), .ZN(n6659) );
  OAI21_X4 U4580 ( .B1(n6752), .B2(n6751), .A(n6750), .ZN(n6753) );
  NAND2_X4 U4581 ( .A1(n4051), .A2(net242080), .ZN(n4035) );
  XNOR2_X1 U4582 ( .A(n8177), .B(n8172), .ZN(n8495) );
  INV_X2 U4583 ( .A(net242079), .ZN(n4052) );
  INV_X8 U4584 ( .A(net242068), .ZN(net241772) );
  INV_X2 U4585 ( .A(n6744), .ZN(n4435) );
  INV_X2 U4586 ( .A(net240930), .ZN(net240939) );
  NAND2_X4 U4587 ( .A1(n4272), .A2(net240951), .ZN(net240933) );
  OAI21_X2 U4588 ( .B1(n3888), .B2(net241014), .A(net241013), .ZN(n4276) );
  INV_X2 U4589 ( .A(n5888), .ZN(n4420) );
  OAI21_X4 U4590 ( .B1(net246357), .B2(net246358), .A(net246359), .ZN(n4015)
         );
  OAI21_X2 U4591 ( .B1(net246357), .B2(net246358), .A(net246359), .ZN(
        net246246) );
  AOI211_X2 U4592 ( .C1(net245893), .C2(net248357), .A(net245895), .B(
        net245896), .ZN(net245892) );
  NOR2_X2 U4593 ( .A1(net245703), .A2(n4073), .ZN(net245697) );
  NOR2_X2 U4594 ( .A1(n5941), .A2(n5083), .ZN(n5943) );
  XNOR2_X2 U4595 ( .A(net246106), .B(net246107), .ZN(n4016) );
  XNOR2_X2 U4596 ( .A(net249297), .B(n4342), .ZN(n4017) );
  XNOR2_X2 U4597 ( .A(n4038), .B(n4219), .ZN(net249297) );
  XNOR2_X2 U4598 ( .A(n7216), .B(n7215), .ZN(n4018) );
  OAI21_X2 U4599 ( .B1(net245994), .B2(net248132), .A(net245897), .ZN(
        net245958) );
  NAND2_X4 U4600 ( .A1(net248132), .A2(net245897), .ZN(net245774) );
  CLKBUF_X3 U4601 ( .A(n7857), .Z(n4027) );
  INV_X1 U4602 ( .A(net246003), .ZN(n4112) );
  XNOR2_X1 U4603 ( .A(n4240), .B(n4241), .ZN(n4019) );
  XNOR2_X2 U4604 ( .A(n4405), .B(n6039), .ZN(n4020) );
  INV_X4 U4605 ( .A(n4020), .ZN(n6086) );
  NAND2_X4 U4606 ( .A1(a[25]), .A2(b[30]), .ZN(n4021) );
  CLKBUF_X3 U4607 ( .A(net245422), .Z(n4022) );
  XNOR2_X1 U4608 ( .A(n6653), .B(n6805), .ZN(n4023) );
  NOR2_X2 U4609 ( .A1(n8456), .A2(n8455), .ZN(n8459) );
  OAI21_X2 U4610 ( .B1(n8521), .B2(n8520), .A(n8519), .ZN(n8523) );
  NAND2_X4 U4611 ( .A1(n7285), .A2(n4382), .ZN(n7596) );
  INV_X4 U4612 ( .A(n7215), .ZN(n4382) );
  OAI22_X4 U4613 ( .A1(net242597), .A2(n7440), .B1(net242602), .B2(n7437), 
        .ZN(n7391) );
  INV_X8 U4614 ( .A(n4103), .ZN(n7387) );
  OAI21_X2 U4615 ( .B1(net240983), .B2(net240961), .A(net240960), .ZN(
        net240980) );
  XNOR2_X2 U4616 ( .A(n4273), .B(net240956), .ZN(n4024) );
  XNOR2_X2 U4617 ( .A(net241586), .B(net241587), .ZN(n4025) );
  AOI21_X4 U4618 ( .B1(net241579), .B2(net242103), .A(n3888), .ZN(n4026) );
  XNOR2_X2 U4619 ( .A(n8096), .B(n7814), .ZN(n4028) );
  XNOR2_X2 U4620 ( .A(n3981), .B(n8150), .ZN(n4029) );
  NAND2_X2 U4621 ( .A1(net242101), .A2(net242102), .ZN(net242366) );
  XNOR2_X2 U4622 ( .A(net241581), .B(net241044), .ZN(n4030) );
  INV_X2 U4623 ( .A(n4124), .ZN(n4031) );
  INV_X4 U4624 ( .A(net240983), .ZN(n4032) );
  NAND2_X4 U4625 ( .A1(net246481), .A2(net246483), .ZN(net246485) );
  NAND2_X4 U4626 ( .A1(b[22]), .A2(net246768), .ZN(net245679) );
  INV_X1 U4627 ( .A(n4034), .ZN(n4033) );
  INV_X1 U4628 ( .A(n4191), .ZN(n4034) );
  OAI21_X2 U4629 ( .B1(net241042), .B2(net249316), .A(n4035), .ZN(net241040)
         );
  NAND2_X4 U4630 ( .A1(net241020), .A2(n4035), .ZN(n4279) );
  NOR2_X4 U4631 ( .A1(net246111), .A2(net246110), .ZN(n4036) );
  INV_X4 U4632 ( .A(net246109), .ZN(net246110) );
  INV_X4 U4633 ( .A(net246475), .ZN(net246470) );
  NAND2_X4 U4634 ( .A1(a[19]), .A2(b[22]), .ZN(n6833) );
  INV_X2 U4635 ( .A(n6087), .ZN(n5925) );
  NOR2_X2 U4636 ( .A1(n6960), .A2(n6959), .ZN(n6963) );
  INV_X2 U4637 ( .A(n6533), .ZN(n6386) );
  NAND2_X2 U4638 ( .A1(n4222), .A2(net245907), .ZN(net245785) );
  OAI22_X2 U4639 ( .A1(net248030), .A2(net248029), .B1(net244274), .B2(
        net244273), .ZN(n4037) );
  AOI22_X2 U4640 ( .A1(net244274), .A2(net244273), .B1(net244553), .B2(
        net244554), .ZN(net244465) );
  INV_X4 U4641 ( .A(net244274), .ZN(net248030) );
  NAND2_X1 U4642 ( .A1(net246760), .A2(b[20]), .ZN(net244554) );
  NAND2_X4 U4643 ( .A1(b[23]), .A2(net246768), .ZN(net245759) );
  XNOR2_X2 U4644 ( .A(n8347), .B(n8562), .ZN(n8756) );
  INV_X2 U4645 ( .A(n8347), .ZN(n8755) );
  NAND2_X4 U4646 ( .A1(n8561), .A2(n8560), .ZN(n8347) );
  INV_X4 U4647 ( .A(n7708), .ZN(n7594) );
  INV_X2 U4648 ( .A(net245744), .ZN(net247658) );
  INV_X1 U4649 ( .A(n7816), .ZN(n7817) );
  XNOR2_X2 U4650 ( .A(n4110), .B(n4090), .ZN(n4038) );
  NOR2_X2 U4651 ( .A1(net242818), .A2(n4217), .ZN(net242821) );
  NAND2_X2 U4652 ( .A1(n7064), .A2(n7063), .ZN(n7072) );
  NAND2_X4 U4653 ( .A1(net243171), .A2(net242894), .ZN(net243167) );
  INV_X2 U4654 ( .A(net243400), .ZN(net243406) );
  INV_X4 U4655 ( .A(net243315), .ZN(net243314) );
  INV_X1 U4656 ( .A(n8279), .ZN(n8276) );
  OAI21_X2 U4657 ( .B1(n4172), .B2(n4017), .A(n4173), .ZN(n4039) );
  NAND2_X2 U4658 ( .A1(net242825), .A2(n4039), .ZN(net242595) );
  INV_X4 U4659 ( .A(net241830), .ZN(net242067) );
  NAND2_X4 U4660 ( .A1(a[28]), .A2(b[10]), .ZN(net242837) );
  INV_X4 U4661 ( .A(n6535), .ZN(n6532) );
  NAND2_X4 U4662 ( .A1(n7620), .A2(net242402), .ZN(n7273) );
  NAND2_X4 U4663 ( .A1(b[19]), .A2(a[24]), .ZN(net243734) );
  AND2_X2 U4664 ( .A1(n7609), .A2(n7608), .ZN(n4040) );
  INV_X4 U4665 ( .A(n4040), .ZN(n7617) );
  NAND2_X2 U4666 ( .A1(n7312), .A2(n7311), .ZN(n7193) );
  NAND2_X4 U4667 ( .A1(n7626), .A2(n7627), .ZN(n7700) );
  NAND2_X4 U4668 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  NOR2_X2 U4669 ( .A1(n4041), .A2(net243639), .ZN(net243637) );
  NOR2_X4 U4670 ( .A1(net243283), .A2(net243284), .ZN(n6938) );
  OAI211_X4 U4671 ( .C1(net242904), .C2(n4219), .A(net242906), .B(net242907), 
        .ZN(net242402) );
  INV_X8 U4672 ( .A(net242909), .ZN(n4219) );
  AOI21_X4 U4673 ( .B1(n6679), .B2(n6680), .A(n6683), .ZN(n4041) );
  INV_X4 U4674 ( .A(n4041), .ZN(n6684) );
  NAND2_X4 U4675 ( .A1(n4052), .A2(n3943), .ZN(n4051) );
  NAND2_X1 U4676 ( .A1(net242100), .A2(n3896), .ZN(n4042) );
  NAND2_X4 U4677 ( .A1(net242100), .A2(net242101), .ZN(net241614) );
  INV_X4 U4678 ( .A(net249128), .ZN(net243433) );
  OAI21_X2 U4679 ( .B1(net241048), .B2(net240997), .A(net240995), .ZN(
        net241047) );
  NOR2_X4 U4680 ( .A1(net243866), .A2(n4292), .ZN(n4290) );
  INV_X8 U4681 ( .A(net243868), .ZN(net243866) );
  NAND2_X2 U4682 ( .A1(n5946), .A2(n5945), .ZN(n6097) );
  INV_X4 U4683 ( .A(n5945), .ZN(n5948) );
  NAND2_X4 U4684 ( .A1(b[15]), .A2(net246766), .ZN(net243401) );
  NAND2_X4 U4685 ( .A1(net241493), .A2(n4158), .ZN(net241593) );
  INV_X4 U4686 ( .A(net243760), .ZN(net243755) );
  NAND2_X4 U4687 ( .A1(b[17]), .A2(net246766), .ZN(net243760) );
  NAND2_X4 U4688 ( .A1(net247549), .A2(n5082), .ZN(n5940) );
  OAI211_X2 U4689 ( .C1(net243866), .C2(net243760), .A(net243761), .B(
        net243757), .ZN(n4043) );
  OAI21_X4 U4690 ( .B1(net242604), .B2(net242603), .A(net242605), .ZN(n4044)
         );
  NOR2_X1 U4691 ( .A1(n7557), .A2(n7556), .ZN(n7560) );
  NAND2_X1 U4692 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  INV_X1 U4693 ( .A(n4307), .ZN(n4046) );
  OAI21_X4 U4694 ( .B1(n6894), .B2(n6893), .A(n6892), .ZN(n4045) );
  NAND2_X2 U4695 ( .A1(n4306), .A2(n4046), .ZN(net242916) );
  XNOR2_X2 U4696 ( .A(n4048), .B(n4047), .ZN(n7538) );
  XNOR2_X2 U4697 ( .A(n7527), .B(n7528), .ZN(n4048) );
  NAND2_X4 U4698 ( .A1(a[24]), .A2(b[16]), .ZN(net243270) );
  INV_X1 U4699 ( .A(n4470), .ZN(n4384) );
  NAND2_X1 U4700 ( .A1(n4307), .A2(net243310), .ZN(net243307) );
  XNOR2_X2 U4701 ( .A(net243175), .B(net243176), .ZN(net248775) );
  XNOR2_X2 U4702 ( .A(n4050), .B(n4049), .ZN(n7967) );
  XNOR2_X2 U4703 ( .A(n7956), .B(n7957), .ZN(n4050) );
  AOI21_X4 U4704 ( .B1(n8539), .B2(n8538), .A(n8540), .ZN(n8162) );
  NOR2_X2 U4705 ( .A1(n3950), .A2(n5958), .ZN(n5962) );
  NOR2_X2 U4706 ( .A1(n3950), .A2(n5959), .ZN(n5956) );
  NAND2_X1 U4707 ( .A1(net243375), .A2(net243376), .ZN(net243186) );
  INV_X4 U4708 ( .A(n6755), .ZN(n6734) );
  INV_X8 U4709 ( .A(net241609), .ZN(net241615) );
  NAND2_X4 U4710 ( .A1(net246772), .A2(b[7]), .ZN(net241609) );
  NAND2_X4 U4711 ( .A1(n4051), .A2(net242080), .ZN(net241021) );
  NAND2_X1 U4712 ( .A1(b[18]), .A2(net246788), .ZN(n5947) );
  OAI21_X2 U4713 ( .B1(net243637), .B2(n4075), .A(net243580), .ZN(net243636)
         );
  INV_X8 U4714 ( .A(net240934), .ZN(n4270) );
  INV_X4 U4715 ( .A(n4933), .ZN(n4931) );
  INV_X4 U4716 ( .A(net241597), .ZN(n4129) );
  NAND2_X1 U4717 ( .A1(n7471), .A2(n7470), .ZN(n7472) );
  XOR2_X1 U4718 ( .A(net241772), .B(net241773), .Z(net249316) );
  NOR2_X4 U4719 ( .A1(net240986), .A2(net241562), .ZN(n4054) );
  INV_X4 U4720 ( .A(n4054), .ZN(net240960) );
  NAND2_X1 U4721 ( .A1(net241568), .A2(net241567), .ZN(net240986) );
  INV_X4 U4722 ( .A(net240985), .ZN(net241562) );
  NAND2_X2 U4723 ( .A1(net241771), .A2(net241770), .ZN(net241045) );
  NAND2_X2 U4724 ( .A1(n6179), .A2(n6178), .ZN(n6070) );
  INV_X1 U4725 ( .A(net240996), .ZN(net241048) );
  XNOR2_X2 U4726 ( .A(n4056), .B(n4055), .ZN(n8406) );
  XNOR2_X2 U4727 ( .A(n8395), .B(n8396), .ZN(n4056) );
  XNOR2_X2 U4728 ( .A(net241817), .B(n4030), .ZN(n4057) );
  XNOR2_X2 U4729 ( .A(n6596), .B(n6544), .ZN(n4436) );
  INV_X2 U4730 ( .A(net240965), .ZN(net241000) );
  NAND2_X4 U4731 ( .A1(net240964), .A2(net240965), .ZN(net240988) );
  XNOR2_X2 U4732 ( .A(n4377), .B(n6257), .ZN(n4434) );
  INV_X4 U4733 ( .A(n6302), .ZN(n4377) );
  INV_X4 U4734 ( .A(n7301), .ZN(n7103) );
  INV_X2 U4735 ( .A(net241014), .ZN(net241010) );
  INV_X2 U4736 ( .A(n8273), .ZN(n8275) );
  NOR2_X2 U4737 ( .A1(n4025), .A2(net241071), .ZN(n4067) );
  NOR2_X2 U4738 ( .A1(n4025), .A2(net241070), .ZN(n4068) );
  NOR2_X4 U4739 ( .A1(n8274), .A2(net241579), .ZN(n7859) );
  INV_X1 U4740 ( .A(net241045), .ZN(net241042) );
  OAI21_X4 U4741 ( .B1(n4027), .B2(n7856), .A(n7855), .ZN(n8273) );
  NAND2_X4 U4742 ( .A1(n4346), .A2(n4347), .ZN(net241020) );
  NAND2_X4 U4743 ( .A1(a[28]), .A2(b[7]), .ZN(net241613) );
  INV_X4 U4744 ( .A(net241071), .ZN(n4058) );
  INV_X1 U4745 ( .A(net241070), .ZN(n4059) );
  NOR2_X2 U4746 ( .A1(n4059), .A2(n4061), .ZN(n4060) );
  NOR2_X2 U4747 ( .A1(n3902), .A2(n3944), .ZN(n4064) );
  NOR2_X4 U4748 ( .A1(n4059), .A2(n4066), .ZN(n4065) );
  NOR2_X4 U4749 ( .A1(n3902), .A2(n4058), .ZN(n4069) );
  INV_X4 U4750 ( .A(n4069), .ZN(n4066) );
  NOR2_X2 U4751 ( .A1(n4064), .A2(n4065), .ZN(n4071) );
  NAND2_X4 U4752 ( .A1(n4070), .A2(n4071), .ZN(n4072) );
  INV_X8 U4753 ( .A(n4072), .ZN(net241022) );
  OAI21_X2 U4754 ( .B1(net245700), .B2(net249328), .A(net245702), .ZN(n5087)
         );
  INV_X2 U4755 ( .A(n4073), .ZN(net245702) );
  OAI21_X1 U4756 ( .B1(n4229), .B2(net249076), .A(net246100), .ZN(n4227) );
  INV_X4 U4757 ( .A(net246446), .ZN(net248353) );
  NAND2_X1 U4758 ( .A1(n7612), .A2(n7611), .ZN(n7613) );
  OAI22_X4 U4759 ( .A1(n7609), .A2(n7608), .B1(n7612), .B2(n7611), .ZN(n7384)
         );
  NOR2_X4 U4760 ( .A1(net245688), .A2(n4170), .ZN(n4164) );
  NOR2_X4 U4761 ( .A1(n5085), .A2(n5084), .ZN(n4073) );
  NAND2_X4 U4762 ( .A1(a[28]), .A2(b[20]), .ZN(n5086) );
  NAND2_X2 U4763 ( .A1(n4677), .A2(n4116), .ZN(n4074) );
  INV_X4 U4764 ( .A(n4074), .ZN(net246570) );
  NAND2_X2 U4765 ( .A1(n7302), .A2(n4408), .ZN(n7303) );
  INV_X4 U4766 ( .A(n4075), .ZN(net243584) );
  NAND2_X4 U4767 ( .A1(a[28]), .A2(b[14]), .ZN(n6683) );
  NAND2_X4 U4768 ( .A1(a[28]), .A2(b[22]), .ZN(net245962) );
  CLKBUF_X2 U4769 ( .A(n5074), .Z(n4459) );
  NOR2_X2 U4770 ( .A1(n7274), .A2(n4076), .ZN(n4096) );
  XNOR2_X2 U4771 ( .A(n7216), .B(n7215), .ZN(n4076) );
  NAND2_X4 U4772 ( .A1(n8260), .A2(n8259), .ZN(n8262) );
  INV_X1 U4773 ( .A(net248549), .ZN(net245209) );
  OAI21_X4 U4774 ( .B1(n4205), .B2(net249300), .A(n4206), .ZN(n4204) );
  NAND2_X4 U4775 ( .A1(n4343), .A2(net243118), .ZN(n4342) );
  INV_X4 U4776 ( .A(net248988), .ZN(net243625) );
  XNOR2_X2 U4777 ( .A(n4078), .B(n4077), .ZN(n7165) );
  XNOR2_X2 U4778 ( .A(n7154), .B(n7155), .ZN(n4078) );
  INV_X8 U4779 ( .A(n6465), .ZN(n6467) );
  XNOR2_X2 U4780 ( .A(n4080), .B(n4079), .ZN(n8366) );
  XNOR2_X2 U4781 ( .A(n8355), .B(n8356), .ZN(n4080) );
  INV_X2 U4782 ( .A(n4081), .ZN(net245616) );
  NAND2_X4 U4783 ( .A1(net244698), .A2(net244697), .ZN(n4082) );
  NAND2_X1 U4784 ( .A1(net244694), .A2(net244695), .ZN(n4083) );
  NAND2_X2 U4785 ( .A1(n4082), .A2(n4083), .ZN(n4081) );
  XNOR2_X2 U4786 ( .A(n4081), .B(n4084), .ZN(net244679) );
  INV_X4 U4787 ( .A(net247491), .ZN(n4084) );
  INV_X8 U4788 ( .A(net245694), .ZN(n4168) );
  NAND2_X2 U4789 ( .A1(b[30]), .A2(a[30]), .ZN(net246579) );
  NAND2_X2 U4790 ( .A1(n4784), .A2(n4376), .ZN(n4712) );
  NAND2_X4 U4791 ( .A1(b[24]), .A2(net246772), .ZN(net245898) );
  INV_X2 U4792 ( .A(net246569), .ZN(n4335) );
  NAND4_X2 U4793 ( .A1(net247667), .A2(b[31]), .A3(a[30]), .A4(a[31]), .ZN(
        n4086) );
  INV_X16 U4794 ( .A(a[29]), .ZN(net247667) );
  NAND2_X1 U4795 ( .A1(b[11]), .A2(net246788), .ZN(net243362) );
  INV_X4 U4796 ( .A(net243313), .ZN(net243361) );
  XNOR2_X2 U4797 ( .A(n7370), .B(n4087), .ZN(n7600) );
  XNOR2_X2 U4798 ( .A(n4089), .B(n4088), .ZN(n7903) );
  XNOR2_X2 U4799 ( .A(n7996), .B(n7999), .ZN(n4089) );
  INV_X2 U4800 ( .A(n6090), .ZN(n6091) );
  NAND2_X4 U4801 ( .A1(b[12]), .A2(a[28]), .ZN(net243181) );
  XNOR2_X2 U4802 ( .A(n4110), .B(n4090), .ZN(net243187) );
  NOR2_X4 U4803 ( .A1(net242835), .A2(net242838), .ZN(net242831) );
  NAND2_X4 U4804 ( .A1(net248038), .A2(n4174), .ZN(n4477) );
  NAND2_X4 U4805 ( .A1(b[9]), .A2(net246766), .ZN(net241760) );
  NOR2_X2 U4806 ( .A1(n4091), .A2(n3908), .ZN(n4092) );
  NOR2_X2 U4807 ( .A1(n7280), .A2(n3945), .ZN(n4093) );
  NOR2_X2 U4808 ( .A1(n4091), .A2(n4100), .ZN(n4095) );
  NOR2_X2 U4809 ( .A1(n4092), .A2(n4093), .ZN(n4097) );
  NOR2_X2 U4810 ( .A1(n4094), .A2(n4095), .ZN(n4098) );
  NAND2_X4 U4811 ( .A1(n4097), .A2(n4098), .ZN(n4099) );
  AND2_X2 U4812 ( .A1(n7223), .A2(n4096), .ZN(n4094) );
  NAND2_X1 U4813 ( .A1(n7223), .A2(n4018), .ZN(n4100) );
  INV_X2 U4814 ( .A(n4018), .ZN(n7280) );
  XNOR2_X2 U4815 ( .A(n4102), .B(n7919), .ZN(n4101) );
  XNOR2_X2 U4816 ( .A(n7916), .B(n7917), .ZN(n4102) );
  XNOR2_X2 U4817 ( .A(n7386), .B(n7385), .ZN(n4103) );
  OAI21_X2 U4818 ( .B1(n7685), .B2(n7684), .A(n3951), .ZN(n7692) );
  AOI21_X2 U4819 ( .B1(n7684), .B2(n3951), .A(n7685), .ZN(n7451) );
  XNOR2_X2 U4820 ( .A(n8279), .B(n8277), .ZN(n8105) );
  NAND2_X4 U4821 ( .A1(n5068), .A2(n5066), .ZN(n4980) );
  NAND2_X4 U4822 ( .A1(n7088), .A2(n7087), .ZN(n7289) );
  NAND2_X4 U4823 ( .A1(n7087), .A2(n7085), .ZN(n7077) );
  NAND2_X4 U4824 ( .A1(n6948), .A2(n6947), .ZN(n7087) );
  INV_X4 U4825 ( .A(net240991), .ZN(net249043) );
  NOR2_X2 U4826 ( .A1(n7114), .A2(n7115), .ZN(n7118) );
  NOR2_X2 U4827 ( .A1(n6824), .A2(n6823), .ZN(n6827) );
  INV_X8 U4828 ( .A(net244379), .ZN(net244153) );
  NAND2_X4 U4829 ( .A1(b[19]), .A2(net246760), .ZN(net244379) );
  INV_X2 U4830 ( .A(net243279), .ZN(net243288) );
  XNOR2_X2 U4831 ( .A(n4398), .B(n4527), .ZN(n4402) );
  INV_X4 U4832 ( .A(net249194), .ZN(net243727) );
  INV_X1 U4833 ( .A(n7362), .ZN(n7366) );
  NAND2_X1 U4834 ( .A1(n6850), .A2(n6851), .ZN(n6852) );
  XNOR2_X2 U4835 ( .A(net240962), .B(net240963), .ZN(n4104) );
  XNOR2_X1 U4836 ( .A(net240953), .B(net240954), .ZN(n4105) );
  NAND2_X4 U4837 ( .A1(n7614), .A2(n7613), .ZN(n7616) );
  INV_X2 U4838 ( .A(n7610), .ZN(n7614) );
  OAI21_X1 U4839 ( .B1(n8579), .B2(n8578), .A(n8577), .ZN(n8738) );
  NOR2_X2 U4840 ( .A1(n7478), .A2(n7477), .ZN(n7481) );
  NAND2_X2 U4841 ( .A1(n7478), .A2(n7477), .ZN(n7479) );
  OAI221_X1 U4842 ( .B1(n5453), .B2(n5452), .C1(net248517), .C2(n5821), .A(
        n5451), .ZN(n5484) );
  NAND2_X1 U4843 ( .A1(n5452), .A2(net246463), .ZN(n4716) );
  XNOR2_X1 U4844 ( .A(n4021), .B(n4767), .ZN(n4700) );
  AOI21_X4 U4845 ( .B1(net245800), .B2(net245801), .A(net245802), .ZN(
        net245794) );
  NOR2_X2 U4846 ( .A1(net245803), .A2(net245804), .ZN(net245800) );
  NAND3_X2 U4847 ( .A1(net243789), .A2(net243790), .A3(net243791), .ZN(n4184)
         );
  NAND2_X2 U4848 ( .A1(net243790), .A2(net243789), .ZN(net243997) );
  NAND2_X4 U4849 ( .A1(n5078), .A2(n5079), .ZN(n5939) );
  INV_X1 U4850 ( .A(n5077), .ZN(n5079) );
  NAND2_X2 U4851 ( .A1(n6875), .A2(n6874), .ZN(n6880) );
  XNOR2_X2 U4852 ( .A(n5009), .B(n4969), .ZN(n5032) );
  INV_X2 U4853 ( .A(n4805), .ZN(n4807) );
  NAND2_X4 U4854 ( .A1(n6038), .A2(n6222), .ZN(n5927) );
  XNOR2_X2 U4855 ( .A(n4772), .B(n4773), .ZN(n4106) );
  INV_X4 U4856 ( .A(n4106), .ZN(n4702) );
  INV_X2 U4857 ( .A(n4772), .ZN(n4785) );
  NAND2_X4 U4858 ( .A1(net245998), .A2(net245898), .ZN(net245997) );
  INV_X1 U4859 ( .A(n6199), .ZN(n6078) );
  AND3_X4 U4860 ( .A1(net246401), .A2(net246402), .A3(net246403), .ZN(n4305)
         );
  NAND2_X4 U4861 ( .A1(n4676), .A2(net246792), .ZN(n4682) );
  INV_X16 U4862 ( .A(net246792), .ZN(net246788) );
  NAND2_X1 U4863 ( .A1(n7371), .A2(n7062), .ZN(n7011) );
  NAND2_X2 U4864 ( .A1(n7129), .A2(n7130), .ZN(n7328) );
  OAI21_X4 U4865 ( .B1(n7128), .B2(n7127), .A(n7126), .ZN(n7130) );
  INV_X4 U4866 ( .A(net240931), .ZN(net240944) );
  NAND2_X2 U4867 ( .A1(net244685), .A2(net245615), .ZN(net245730) );
  NAND2_X4 U4868 ( .A1(net240929), .A2(net240930), .ZN(net240928) );
  INV_X8 U4869 ( .A(net241031), .ZN(n4299) );
  XNOR2_X2 U4870 ( .A(n4318), .B(n3890), .ZN(net243743) );
  NAND2_X4 U4871 ( .A1(n4228), .A2(net246086), .ZN(n4224) );
  NAND2_X4 U4872 ( .A1(n4016), .A2(n4227), .ZN(n4226) );
  OAI21_X4 U4873 ( .B1(n3966), .B2(net245981), .A(n4929), .ZN(n4933) );
  XOR2_X2 U4874 ( .A(net246540), .B(net246506), .Z(net246537) );
  INV_X2 U4875 ( .A(net246016), .ZN(net246014) );
  INV_X4 U4876 ( .A(net245738), .ZN(net248083) );
  NAND2_X4 U4877 ( .A1(net246836), .A2(a[28]), .ZN(net245738) );
  XNOR2_X2 U4878 ( .A(n4105), .B(net240932), .ZN(net240927) );
  AOI21_X2 U4879 ( .B1(net244689), .B2(net244690), .A(n4309), .ZN(net244687)
         );
  NAND2_X2 U4880 ( .A1(n4107), .A2(n4108), .ZN(n4109) );
  INV_X1 U4881 ( .A(n4013), .ZN(n4107) );
  INV_X4 U4882 ( .A(n4109), .ZN(n7188) );
  NAND2_X4 U4883 ( .A1(net242917), .A2(net242916), .ZN(n4110) );
  OAI22_X2 U4884 ( .A1(net246535), .A2(net246534), .B1(net246530), .B2(n4355), 
        .ZN(net246516) );
  INV_X4 U4885 ( .A(n4116), .ZN(net246535) );
  NAND2_X2 U4886 ( .A1(net246110), .A2(net246111), .ZN(net246004) );
  NAND2_X4 U4887 ( .A1(n4830), .A2(net246100), .ZN(net246186) );
  OAI21_X4 U4888 ( .B1(n7800), .B2(n4525), .A(n7799), .ZN(n7441) );
  NAND2_X4 U4889 ( .A1(net240783), .A2(n4358), .ZN(net240925) );
  NAND2_X4 U4890 ( .A1(n7276), .A2(n7275), .ZN(n7223) );
  OAI211_X4 U4891 ( .C1(net246537), .C2(net246536), .A(net245393), .B(
        net246538), .ZN(net246515) );
  INV_X8 U4892 ( .A(net246543), .ZN(net246536) );
  NAND2_X4 U4893 ( .A1(a[25]), .A2(b[31]), .ZN(net246463) );
  NAND2_X2 U4894 ( .A1(n4799), .A2(n4800), .ZN(n4111) );
  INV_X4 U4895 ( .A(n4111), .ZN(net248925) );
  AOI21_X4 U4896 ( .B1(n7796), .B2(n8083), .A(n7795), .ZN(n7797) );
  INV_X4 U4897 ( .A(n8081), .ZN(n7795) );
  OAI21_X2 U4898 ( .B1(n4112), .B2(n4113), .A(net249274), .ZN(n4114) );
  INV_X1 U4899 ( .A(net246004), .ZN(n4113) );
  INV_X4 U4900 ( .A(n4114), .ZN(net246107) );
  XNOR2_X2 U4901 ( .A(n4878), .B(n4016), .ZN(net245985) );
  AOI21_X4 U4902 ( .B1(net246177), .B2(net246176), .A(net245429), .ZN(n4115)
         );
  INV_X4 U4903 ( .A(n4115), .ZN(net246017) );
  NAND4_X4 U4904 ( .A1(net247667), .A2(b[31]), .A3(a[30]), .A4(a[31]), .ZN(
        net246582) );
  NAND2_X4 U4905 ( .A1(b[29]), .A2(a[29]), .ZN(net245313) );
  OAI21_X4 U4906 ( .B1(n4678), .B2(n5266), .A(n5294), .ZN(n4116) );
  XNOR2_X2 U4907 ( .A(net246365), .B(net246361), .ZN(net246392) );
  OAI211_X2 U4908 ( .C1(net241607), .C2(net241606), .A(net241608), .B(
        net241609), .ZN(net241588) );
  NAND3_X2 U4909 ( .A1(net245773), .A2(net245774), .A3(net245775), .ZN(
        net245766) );
  OAI21_X4 U4910 ( .B1(net245672), .B2(net245673), .A(net245674), .ZN(
        net244702) );
  INV_X4 U4911 ( .A(net245675), .ZN(net245672) );
  NOR2_X4 U4912 ( .A1(n5870), .A2(n4439), .ZN(n5884) );
  NOR2_X4 U4913 ( .A1(n4899), .A2(n4898), .ZN(n4901) );
  INV_X4 U4914 ( .A(n4895), .ZN(n4899) );
  OAI21_X4 U4915 ( .B1(n5922), .B2(n5921), .A(n5920), .ZN(n5923) );
  INV_X1 U4916 ( .A(n5918), .ZN(n5922) );
  INV_X8 U4917 ( .A(n5914), .ZN(n5921) );
  INV_X1 U4918 ( .A(n5919), .ZN(n5920) );
  OAI21_X4 U4919 ( .B1(net245901), .B2(net248800), .A(net245902), .ZN(
        net245998) );
  CLKBUF_X3 U4920 ( .A(n4036), .Z(net248800) );
  INV_X8 U4921 ( .A(net246002), .ZN(net245902) );
  AOI21_X2 U4922 ( .B1(net245465), .B2(n4182), .A(n3929), .ZN(n4117) );
  INV_X4 U4923 ( .A(n4117), .ZN(net246482) );
  OAI21_X4 U4924 ( .B1(n6320), .B2(n6319), .A(n6318), .ZN(n6438) );
  NAND2_X2 U4925 ( .A1(a[18]), .A2(n5869), .ZN(n6072) );
  OAI211_X4 U4926 ( .C1(n4951), .C2(n4950), .A(n4948), .B(n4949), .ZN(n5029)
         );
  INV_X1 U4927 ( .A(n4945), .ZN(n4951) );
  OAI21_X2 U4928 ( .B1(net246327), .B2(n4761), .A(n4716), .ZN(n4721) );
  NAND2_X4 U4929 ( .A1(n4912), .A2(net246034), .ZN(n4945) );
  NAND3_X4 U4930 ( .A1(n4118), .A2(n5025), .A3(n5040), .ZN(n5088) );
  INV_X2 U4931 ( .A(n5042), .ZN(n4118) );
  NOR3_X4 U4932 ( .A1(n4718), .A2(net247778), .A3(n4119), .ZN(n4720) );
  INV_X4 U4933 ( .A(net246332), .ZN(n4119) );
  INV_X8 U4934 ( .A(n4717), .ZN(n4718) );
  OAI21_X4 U4935 ( .B1(net246243), .B2(net246244), .A(n3930), .ZN(net246176)
         );
  INV_X4 U4936 ( .A(net246248), .ZN(net246243) );
  XNOR2_X2 U4937 ( .A(n7177), .B(n7175), .ZN(n4120) );
  INV_X4 U4938 ( .A(n4120), .ZN(n7002) );
  NAND2_X4 U4939 ( .A1(net246452), .A2(net248742), .ZN(net246448) );
  NAND2_X2 U4940 ( .A1(n7061), .A2(n7060), .ZN(n4515) );
  NAND3_X2 U4941 ( .A1(net246450), .A2(a[29]), .A3(b[28]), .ZN(net246518) );
  NAND2_X2 U4942 ( .A1(net245911), .A2(net245910), .ZN(net245909) );
  OAI21_X2 U4943 ( .B1(n4121), .B2(n4899), .A(n4900), .ZN(n4122) );
  INV_X1 U4944 ( .A(n4858), .ZN(n4121) );
  INV_X2 U4945 ( .A(n4122), .ZN(n4888) );
  OAI21_X4 U4946 ( .B1(n7074), .B2(n4419), .A(n7371), .ZN(n7075) );
  NAND2_X4 U4947 ( .A1(n4336), .A2(n4337), .ZN(net246559) );
  XNOR2_X2 U4948 ( .A(n4684), .B(n4692), .ZN(net246446) );
  XNOR2_X2 U4949 ( .A(n4726), .B(n4756), .ZN(n4729) );
  OAI21_X4 U4950 ( .B1(net246804), .B2(n4123), .A(a[29]), .ZN(net246581) );
  INV_X8 U4951 ( .A(b[31]), .ZN(n4123) );
  NAND3_X2 U4952 ( .A1(net245785), .A2(net245786), .A3(n4124), .ZN(n4125) );
  INV_X4 U4953 ( .A(n4125), .ZN(n5060) );
  OAI21_X4 U4954 ( .B1(net243769), .B2(n4183), .A(net243770), .ZN(net243423)
         );
  INV_X1 U4955 ( .A(net243863), .ZN(n4183) );
  INV_X32 U4956 ( .A(b[3]), .ZN(n8281) );
  OAI21_X4 U4957 ( .B1(n6589), .B2(n6590), .A(n6588), .ZN(net243376) );
  AOI22_X4 U4958 ( .A1(net243295), .A2(net243297), .B1(net243580), .B2(
        net243300), .ZN(net243579) );
  NAND2_X1 U4959 ( .A1(net244275), .A2(net244465), .ZN(net247927) );
  NAND2_X4 U4960 ( .A1(net241068), .A2(net241067), .ZN(net241586) );
  OAI22_X2 U4961 ( .A1(net242069), .A2(net241609), .B1(net241616), .B2(
        net241615), .ZN(net242068) );
  NAND2_X1 U4962 ( .A1(net241615), .A2(net241616), .ZN(net247473) );
  NAND2_X4 U4963 ( .A1(net241588), .A2(net241589), .ZN(net241068) );
  XNOR2_X2 U4964 ( .A(n4126), .B(n4127), .ZN(net241589) );
  XNOR2_X2 U4965 ( .A(n4128), .B(net241593), .ZN(n4127) );
  NAND3_X2 U4966 ( .A1(net241594), .A2(net241595), .A3(net241596), .ZN(n4128)
         );
  NAND2_X4 U4967 ( .A1(n4130), .A2(n4131), .ZN(n4126) );
  NAND2_X4 U4968 ( .A1(net247912), .A2(n4129), .ZN(n4131) );
  INV_X4 U4969 ( .A(net241598), .ZN(net247912) );
  NAND2_X2 U4970 ( .A1(net241598), .A2(net241597), .ZN(n4130) );
  NOR2_X4 U4971 ( .A1(net241610), .A2(net241611), .ZN(net241606) );
  NAND2_X2 U4972 ( .A1(net241612), .A2(net241613), .ZN(net241611) );
  OAI21_X4 U4973 ( .B1(net242070), .B2(net241607), .A(net241608), .ZN(
        net241616) );
  INV_X4 U4974 ( .A(net242077), .ZN(net242070) );
  NAND3_X2 U4975 ( .A1(net241612), .A2(net241614), .A3(net241613), .ZN(
        net242077) );
  INV_X32 U4976 ( .A(net246776), .ZN(net246772) );
  INV_X32 U4977 ( .A(a[27]), .ZN(net246776) );
  XOR2_X2 U4978 ( .A(net241492), .B(net241593), .Z(net241751) );
  NAND3_X2 U4979 ( .A1(net241595), .A2(net241596), .A3(net241594), .ZN(
        net241821) );
  NAND2_X4 U4980 ( .A1(net241614), .A2(net241612), .ZN(net242072) );
  NAND2_X4 U4981 ( .A1(net246399), .A2(net246398), .ZN(net246476) );
  XNOR2_X2 U4982 ( .A(net246476), .B(net246400), .ZN(net246439) );
  NAND2_X4 U4983 ( .A1(net246477), .A2(net246478), .ZN(net246399) );
  NAND2_X1 U4984 ( .A1(net246399), .A2(net246398), .ZN(net246395) );
  OAI21_X4 U4985 ( .B1(net246479), .B2(net246480), .A(net246481), .ZN(
        net246478) );
  INV_X4 U4986 ( .A(net246482), .ZN(net246480) );
  INV_X4 U4987 ( .A(net246491), .ZN(net246479) );
  NAND2_X1 U4988 ( .A1(net248913), .A2(net246479), .ZN(net247815) );
  INV_X1 U4989 ( .A(net246479), .ZN(net249130) );
  NOR2_X4 U4990 ( .A1(net246479), .A2(net246488), .ZN(net246484) );
  INV_X4 U4991 ( .A(net246483), .ZN(net246477) );
  OAI21_X4 U4992 ( .B1(net246484), .B2(net246485), .A(net246486), .ZN(
        net246398) );
  INV_X4 U4993 ( .A(net246487), .ZN(net246486) );
  INV_X1 U4994 ( .A(net246486), .ZN(net249142) );
  XNOR2_X2 U4995 ( .A(net246502), .B(n4132), .ZN(net246487) );
  NAND3_X2 U4996 ( .A1(net246518), .A2(net246448), .A3(n4133), .ZN(n4132) );
  NAND2_X1 U4997 ( .A1(net246450), .A2(net248742), .ZN(n4133) );
  INV_X8 U4998 ( .A(net246522), .ZN(net246450) );
  XNOR2_X2 U4999 ( .A(net246468), .B(n4134), .ZN(net246522) );
  XNOR2_X2 U5000 ( .A(n4135), .B(n4136), .ZN(n4134) );
  INV_X4 U5001 ( .A(net246516), .ZN(n4136) );
  NAND2_X2 U5002 ( .A1(net247797), .A2(n4137), .ZN(n4135) );
  NAND2_X2 U5003 ( .A1(net247795), .A2(net248379), .ZN(n4137) );
  INV_X4 U5004 ( .A(net245349), .ZN(net246467) );
  NAND2_X2 U5005 ( .A1(net246467), .A2(net246468), .ZN(net246466) );
  NAND2_X4 U5006 ( .A1(net246468), .A2(net246467), .ZN(net246475) );
  NAND2_X2 U5007 ( .A1(net246467), .A2(net246517), .ZN(net247797) );
  INV_X4 U5008 ( .A(net248379), .ZN(net246517) );
  XNOR2_X2 U5009 ( .A(net246516), .B(net246517), .ZN(net246511) );
  NAND2_X4 U5010 ( .A1(net245958), .A2(net245893), .ZN(net245957) );
  XNOR2_X2 U5011 ( .A(net245957), .B(net245773), .ZN(net245956) );
  NAND2_X1 U5012 ( .A1(net245893), .A2(net245958), .ZN(net245993) );
  INV_X4 U5013 ( .A(net245997), .ZN(net245994) );
  NAND3_X2 U5014 ( .A1(net245766), .A2(net245893), .A3(net247540), .ZN(
        net245768) );
  NAND2_X2 U5015 ( .A1(net245766), .A2(net245893), .ZN(net245765) );
  NOR2_X4 U5016 ( .A1(net248132), .A2(net245897), .ZN(net245904) );
  NAND3_X2 U5017 ( .A1(net245897), .A2(net245898), .A3(net245899), .ZN(
        net245775) );
  NAND2_X2 U5018 ( .A1(net245898), .A2(net245998), .ZN(net245905) );
  XNOR2_X2 U5019 ( .A(net245902), .B(net245898), .ZN(net246106) );
  NAND2_X4 U5020 ( .A1(net246520), .A2(net246521), .ZN(net247186) );
  XNOR2_X2 U5021 ( .A(net247186), .B(net246523), .ZN(net246526) );
  NAND2_X2 U5022 ( .A1(net246549), .A2(net247173), .ZN(net246520) );
  NAND2_X4 U5023 ( .A1(net246520), .A2(net246521), .ZN(net248742) );
  OAI21_X4 U5024 ( .B1(net247173), .B2(net246549), .A(net246550), .ZN(
        net246521) );
  XNOR2_X2 U5025 ( .A(net246560), .B(net246559), .ZN(net246550) );
  INV_X4 U5026 ( .A(net246551), .ZN(net246549) );
  XNOR2_X2 U5027 ( .A(net247173), .B(net246551), .ZN(net246557) );
  XNOR2_X1 U5028 ( .A(net246560), .B(net246559), .ZN(net248717) );
  NAND2_X4 U5029 ( .A1(net240964), .A2(net240965), .ZN(net240963) );
  XNOR2_X2 U5030 ( .A(net240962), .B(net240963), .ZN(net240953) );
  NAND2_X2 U5031 ( .A1(net241001), .A2(net241002), .ZN(net240964) );
  OAI21_X2 U5032 ( .B1(net248695), .B2(net241000), .A(net240964), .ZN(
        net240999) );
  INV_X4 U5033 ( .A(net241003), .ZN(net241001) );
  NAND2_X4 U5034 ( .A1(net241004), .A2(net241003), .ZN(net240965) );
  INV_X4 U5035 ( .A(net241002), .ZN(net241004) );
  INV_X4 U5036 ( .A(net242325), .ZN(net242100) );
  OAI21_X2 U5037 ( .B1(net242099), .B2(net242100), .A(n3896), .ZN(net242098)
         );
  XNOR2_X2 U5038 ( .A(net242375), .B(net242376), .ZN(net242325) );
  NAND2_X4 U5039 ( .A1(net242368), .A2(net242367), .ZN(net242101) );
  INV_X2 U5040 ( .A(net242324), .ZN(net242368) );
  XNOR2_X2 U5041 ( .A(net242382), .B(net242314), .ZN(net242375) );
  XNOR2_X1 U5042 ( .A(net242375), .B(net242376), .ZN(net248078) );
  XNOR2_X2 U5043 ( .A(net242383), .B(net242304), .ZN(net242382) );
  AOI22_X2 U5044 ( .A1(net242320), .A2(net242321), .B1(net242303), .B2(
        net242302), .ZN(net242383) );
  INV_X4 U5045 ( .A(net242321), .ZN(net242302) );
  NAND2_X2 U5046 ( .A1(net242302), .A2(net242303), .ZN(net241830) );
  INV_X8 U5047 ( .A(n4044), .ZN(net242320) );
  AND2_X2 U5048 ( .A1(net242320), .A2(net242321), .ZN(net248788) );
  NOR2_X1 U5049 ( .A1(net242320), .A2(net242321), .ZN(net242319) );
  INV_X8 U5050 ( .A(net242377), .ZN(n4138) );
  NOR2_X4 U5051 ( .A1(n4138), .A2(net242315), .ZN(net242309) );
  OAI21_X4 U5052 ( .B1(n4138), .B2(net242311), .A(net242313), .ZN(net242310)
         );
  OAI21_X4 U5053 ( .B1(net242378), .B2(net242379), .A(n4139), .ZN(net242377)
         );
  INV_X4 U5054 ( .A(n4140), .ZN(n4139) );
  INV_X4 U5055 ( .A(n4139), .ZN(net248749) );
  XNOR2_X2 U5056 ( .A(net242666), .B(net242667), .ZN(n4140) );
  NAND2_X1 U5057 ( .A1(net249292), .A2(net242610), .ZN(net242667) );
  INV_X1 U5058 ( .A(net242607), .ZN(net249292) );
  INV_X8 U5059 ( .A(net242613), .ZN(net242607) );
  NOR2_X4 U5060 ( .A1(net246241), .A2(n3852), .ZN(n4141) );
  XNOR2_X2 U5061 ( .A(n4141), .B(n3930), .ZN(net246277) );
  NOR2_X4 U5062 ( .A1(net246242), .A2(net246241), .ZN(net246254) );
  INV_X8 U5063 ( .A(net246247), .ZN(net246241) );
  OAI21_X4 U5064 ( .B1(net246241), .B2(net246242), .A(net246243), .ZN(
        net246177) );
  NAND2_X1 U5065 ( .A1(net246246), .A2(net246247), .ZN(net246244) );
  NAND2_X2 U5066 ( .A1(net246360), .A2(net246361), .ZN(net246358) );
  NAND2_X2 U5067 ( .A1(net246437), .A2(net246436), .ZN(net246360) );
  INV_X4 U5068 ( .A(net246390), .ZN(net246436) );
  NAND2_X2 U5069 ( .A1(net246436), .A2(net246437), .ZN(net247619) );
  NAND2_X4 U5070 ( .A1(net246388), .A2(net246436), .ZN(net246362) );
  NAND2_X4 U5071 ( .A1(net246362), .A2(net246363), .ZN(net246357) );
  NAND2_X4 U5072 ( .A1(net246365), .A2(net246364), .ZN(net246247) );
  INV_X4 U5073 ( .A(net246361), .ZN(net246364) );
  INV_X1 U5074 ( .A(net246359), .ZN(net246393) );
  NAND2_X4 U5075 ( .A1(net246388), .A2(net246437), .ZN(net246363) );
  XNOR2_X2 U5076 ( .A(net246389), .B(net246390), .ZN(net246387) );
  NAND3_X4 U5077 ( .A1(net246363), .A2(net246362), .A3(net247619), .ZN(
        net246365) );
  INV_X4 U5078 ( .A(net246438), .ZN(net246388) );
  INV_X2 U5079 ( .A(net246388), .ZN(net247821) );
  XNOR2_X2 U5080 ( .A(net246439), .B(n4019), .ZN(net246438) );
  NAND2_X2 U5081 ( .A1(net246397), .A2(net246396), .ZN(net246288) );
  NAND2_X2 U5082 ( .A1(net246395), .A2(net246396), .ZN(net246287) );
  INV_X4 U5083 ( .A(net246400), .ZN(net246397) );
  NAND2_X4 U5084 ( .A1(net244383), .A2(net244385), .ZN(net244381) );
  NAND3_X2 U5085 ( .A1(net244380), .A2(net244382), .A3(net244381), .ZN(
        net244154) );
  NAND3_X2 U5086 ( .A1(net244380), .A2(net244382), .A3(net244381), .ZN(
        net247924) );
  INV_X4 U5087 ( .A(net244387), .ZN(net244385) );
  NAND2_X2 U5088 ( .A1(net244384), .A2(net244385), .ZN(net244380) );
  INV_X8 U5089 ( .A(net244386), .ZN(net244383) );
  NAND2_X4 U5090 ( .A1(net244383), .A2(net244384), .ZN(net244382) );
  NAND2_X2 U5091 ( .A1(b[19]), .A2(net246768), .ZN(net244387) );
  XNOR2_X2 U5092 ( .A(net244386), .B(net244387), .ZN(net244457) );
  INV_X8 U5093 ( .A(net246770), .ZN(net246768) );
  INV_X32 U5094 ( .A(a[26]), .ZN(net246770) );
  INV_X32 U5095 ( .A(b[19]), .ZN(n4145) );
  NOR3_X4 U5096 ( .A1(net248549), .A2(net246812), .A3(n4145), .ZN(net245722)
         );
  NAND2_X4 U5097 ( .A1(net247927), .A2(net247928), .ZN(net244386) );
  NAND2_X4 U5098 ( .A1(n4037), .A2(net247926), .ZN(net247928) );
  INV_X4 U5099 ( .A(net244466), .ZN(net244275) );
  NAND2_X2 U5100 ( .A1(net248031), .A2(net244275), .ZN(net244271) );
  XNOR2_X2 U5101 ( .A(n4143), .B(n4142), .ZN(net244466) );
  INV_X4 U5102 ( .A(net244146), .ZN(n4142) );
  NAND3_X2 U5103 ( .A1(n4142), .A2(a[23]), .A3(net244144), .ZN(net244281) );
  XNOR2_X2 U5104 ( .A(net247544), .B(n4144), .ZN(n4143) );
  XNOR2_X2 U5105 ( .A(n4146), .B(net244288), .ZN(n4144) );
  INV_X8 U5106 ( .A(net244372), .ZN(n4146) );
  XNOR2_X2 U5107 ( .A(net244288), .B(n4146), .ZN(net244283) );
  INV_X4 U5108 ( .A(net244289), .ZN(net244372) );
  NOR3_X4 U5109 ( .A1(net240774), .A2(net240775), .A3(n4147), .ZN(zero_signal)
         );
  NAND2_X2 U5110 ( .A1(n4148), .A2(net240767), .ZN(n4147) );
  NOR2_X4 U5111 ( .A1(net240772), .A2(n3952), .ZN(n4148) );
  NAND2_X2 U5112 ( .A1(n4150), .A2(n4151), .ZN(n4149) );
  NAND2_X2 U5113 ( .A1(n4153), .A2(n4154), .ZN(n4152) );
  INV_X4 U5114 ( .A(out[10]), .ZN(n4154) );
  NOR2_X4 U5115 ( .A1(out[11]), .A2(n3971), .ZN(n4153) );
  INV_X4 U5116 ( .A(n4156), .ZN(n4155) );
  NOR2_X4 U5117 ( .A1(out[15]), .A2(n4157), .ZN(n4156) );
  INV_X8 U5118 ( .A(net241746), .ZN(n4158) );
  NAND2_X4 U5119 ( .A1(net241493), .A2(n4158), .ZN(net241832) );
  INV_X1 U5120 ( .A(n4158), .ZN(net241491) );
  NAND2_X4 U5121 ( .A1(n4161), .A2(n4162), .ZN(net241594) );
  NAND2_X2 U5122 ( .A1(n4160), .A2(net241760), .ZN(n4162) );
  INV_X2 U5123 ( .A(net241824), .ZN(n4160) );
  NOR2_X2 U5124 ( .A1(n4160), .A2(n4159), .ZN(net241757) );
  NOR2_X4 U5125 ( .A1(n4159), .A2(net241754), .ZN(n4161) );
  INV_X4 U5126 ( .A(n4028), .ZN(n4159) );
  NOR2_X2 U5127 ( .A1(n4159), .A2(net241760), .ZN(net241758) );
  XNOR2_X2 U5128 ( .A(net242153), .B(n4159), .ZN(net242074) );
  OAI22_X4 U5129 ( .A1(net241749), .A2(net241756), .B1(net241827), .B2(
        net241828), .ZN(net241595) );
  NAND2_X4 U5130 ( .A1(net243746), .A2(net243745), .ZN(net243749) );
  INV_X2 U5131 ( .A(net243749), .ZN(net243747) );
  XNOR2_X2 U5132 ( .A(net243749), .B(net243578), .ZN(net243874) );
  OAI21_X4 U5133 ( .B1(net243993), .B2(net243994), .A(net243995), .ZN(
        net243746) );
  INV_X1 U5134 ( .A(net243746), .ZN(net243740) );
  INV_X4 U5135 ( .A(net244156), .ZN(net243993) );
  NAND2_X2 U5136 ( .A1(net243993), .A2(net243994), .ZN(net243745) );
  OAI22_X2 U5137 ( .A1(net244155), .A2(net244156), .B1(net243994), .B2(
        net243993), .ZN(net244066) );
  NAND2_X1 U5138 ( .A1(net243745), .A2(net243578), .ZN(net243741) );
  INV_X1 U5139 ( .A(net243994), .ZN(net244155) );
  NAND2_X4 U5140 ( .A1(n4163), .A2(net245681), .ZN(net245676) );
  NAND2_X4 U5141 ( .A1(net245676), .A2(net245677), .ZN(net244694) );
  NAND2_X1 U5142 ( .A1(net245677), .A2(net245676), .ZN(net249197) );
  XNOR2_X2 U5143 ( .A(n4166), .B(net248472), .ZN(net245681) );
  OAI22_X2 U5144 ( .A1(n4167), .A2(net245694), .B1(n4168), .B2(net245696), 
        .ZN(n4166) );
  NAND2_X4 U5145 ( .A1(n4168), .A2(net245696), .ZN(net245675) );
  INV_X4 U5146 ( .A(net245696), .ZN(n4167) );
  NAND2_X2 U5147 ( .A1(n4167), .A2(net245694), .ZN(net245674) );
  OAI21_X4 U5148 ( .B1(net245683), .B2(n4164), .A(n4165), .ZN(n4163) );
  INV_X4 U5149 ( .A(net245679), .ZN(n4165) );
  INV_X4 U5150 ( .A(n4169), .ZN(n4170) );
  NOR2_X2 U5151 ( .A1(net245687), .A2(net245686), .ZN(n4169) );
  INV_X4 U5152 ( .A(net245690), .ZN(net245687) );
  INV_X2 U5153 ( .A(net245687), .ZN(net249331) );
  INV_X2 U5154 ( .A(net245689), .ZN(net245688) );
  INV_X4 U5155 ( .A(net245691), .ZN(net245683) );
  XNOR2_X2 U5156 ( .A(net245760), .B(n4171), .ZN(net248472) );
  XNOR2_X1 U5157 ( .A(net248472), .B(net245752), .ZN(net245740) );
  CLKBUF_X3 U5158 ( .A(net245621), .Z(n4171) );
  XNOR2_X2 U5159 ( .A(net245760), .B(n4171), .ZN(net245673) );
  NAND3_X4 U5160 ( .A1(net245754), .A2(net245755), .A3(net245753), .ZN(
        net245694) );
  INV_X4 U5161 ( .A(net245759), .ZN(net245758) );
  NAND2_X2 U5162 ( .A1(net245758), .A2(net245757), .ZN(net245754) );
  NAND2_X2 U5163 ( .A1(net245757), .A2(net245756), .ZN(net245755) );
  NAND2_X2 U5164 ( .A1(b[23]), .A2(net246760), .ZN(net245696) );
  INV_X32 U5165 ( .A(net246762), .ZN(net246760) );
  INV_X32 U5166 ( .A(a[25]), .ZN(net246762) );
  NOR2_X4 U5167 ( .A1(net242607), .A2(net242612), .ZN(net242603) );
  NAND2_X4 U5168 ( .A1(net247915), .A2(net248777), .ZN(net242613) );
  OR2_X2 U5169 ( .A1(net242669), .A2(net242668), .ZN(net247915) );
  INV_X4 U5170 ( .A(net242884), .ZN(net242668) );
  NAND2_X2 U5171 ( .A1(net242668), .A2(net242885), .ZN(net242882) );
  NAND2_X2 U5172 ( .A1(net242668), .A2(net242669), .ZN(net242610) );
  INV_X1 U5173 ( .A(net242610), .ZN(net242606) );
  NAND2_X2 U5174 ( .A1(b[9]), .A2(a[28]), .ZN(net242609) );
  XNOR2_X2 U5175 ( .A(net242611), .B(net242609), .ZN(net242666) );
  INV_X4 U5176 ( .A(net242609), .ZN(net242608) );
  XNOR2_X2 U5177 ( .A(net242891), .B(net248778), .ZN(net248777) );
  INV_X2 U5178 ( .A(net248777), .ZN(net248651) );
  OR2_X1 U5179 ( .A1(net242834), .A2(net242835), .ZN(net248778) );
  INV_X4 U5180 ( .A(net242839), .ZN(net242834) );
  OAI21_X4 U5181 ( .B1(net242835), .B2(net242834), .A(net242836), .ZN(
        net242833) );
  XNOR2_X2 U5182 ( .A(net242832), .B(net242837), .ZN(net242891) );
  INV_X4 U5183 ( .A(net242885), .ZN(net242673) );
  OAI211_X1 U5184 ( .C1(net242672), .C2(net242673), .A(net242674), .B(
        net242884), .ZN(net242883) );
  NAND2_X2 U5185 ( .A1(b[9]), .A2(net246788), .ZN(net242884) );
  INV_X32 U5186 ( .A(a[29]), .ZN(net246792) );
  NAND2_X2 U5187 ( .A1(net242839), .A2(net242837), .ZN(net242838) );
  OAI21_X4 U5188 ( .B1(net242831), .B2(net242832), .A(net242833), .ZN(
        net242602) );
  INV_X4 U5189 ( .A(net242837), .ZN(net242836) );
  XNOR2_X2 U5190 ( .A(net243159), .B(net242672), .ZN(net242879) );
  NOR2_X4 U5191 ( .A1(net243111), .A2(n4175), .ZN(n4172) );
  OAI21_X4 U5192 ( .B1(n4172), .B2(net243108), .A(n4173), .ZN(net242826) );
  NAND2_X2 U5193 ( .A1(net243114), .A2(net243113), .ZN(n4175) );
  INV_X4 U5194 ( .A(net243121), .ZN(net243111) );
  OAI21_X4 U5195 ( .B1(net243111), .B2(net243110), .A(n4174), .ZN(n4173) );
  NAND2_X2 U5196 ( .A1(n4177), .A2(net243313), .ZN(net243114) );
  INV_X4 U5197 ( .A(net243114), .ZN(net243110) );
  NAND2_X4 U5198 ( .A1(net243121), .A2(net243114), .ZN(net243311) );
  INV_X2 U5199 ( .A(net243362), .ZN(n4177) );
  OAI22_X2 U5200 ( .A1(net243361), .A2(net243362), .B1(n4177), .B2(net243313), 
        .ZN(n4178) );
  NAND2_X4 U5201 ( .A1(b[11]), .A2(a[28]), .ZN(net243113) );
  INV_X4 U5202 ( .A(net243113), .ZN(n4174) );
  NAND2_X4 U5203 ( .A1(net243314), .A2(n4179), .ZN(net243121) );
  XNOR2_X2 U5204 ( .A(net243314), .B(n4178), .ZN(net248693) );
  XNOR2_X2 U5205 ( .A(net243369), .B(net243180), .ZN(net243315) );
  INV_X4 U5206 ( .A(net243370), .ZN(net243180) );
  NAND2_X4 U5207 ( .A1(net243180), .A2(net243181), .ZN(net243179) );
  NAND2_X2 U5208 ( .A1(net243186), .A2(net243185), .ZN(net243370) );
  XNOR2_X2 U5209 ( .A(net243377), .B(net243378), .ZN(n4176) );
  XNOR2_X2 U5210 ( .A(net243378), .B(net243377), .ZN(net248703) );
  INV_X4 U5211 ( .A(n4181), .ZN(n4180) );
  NAND2_X4 U5212 ( .A1(n4180), .A2(n3929), .ZN(net246481) );
  XNOR2_X2 U5213 ( .A(n4181), .B(n3929), .ZN(net248913) );
  NAND2_X4 U5214 ( .A1(n4182), .A2(net245465), .ZN(n4181) );
  NOR2_X4 U5215 ( .A1(net247632), .A2(net246874), .ZN(n4182) );
  INV_X32 U5216 ( .A(b[27]), .ZN(net246874) );
  INV_X32 U5217 ( .A(a[31]), .ZN(net247632) );
  XNOR2_X2 U5218 ( .A(net246526), .B(net248571), .ZN(net246491) );
  NAND2_X2 U5219 ( .A1(net246482), .A2(net246491), .ZN(net246497) );
  INV_X2 U5220 ( .A(net246450), .ZN(net248571) );
  NAND2_X4 U5221 ( .A1(net243787), .A2(n4184), .ZN(net243407) );
  NAND2_X2 U5222 ( .A1(net243408), .A2(net243407), .ZN(net243400) );
  NAND2_X4 U5223 ( .A1(net243407), .A2(net243408), .ZN(net243782) );
  INV_X4 U5224 ( .A(net243788), .ZN(net243787) );
  XNOR2_X2 U5225 ( .A(net243861), .B(net243862), .ZN(net243788) );
  XNOR2_X2 U5226 ( .A(net243860), .B(net243788), .ZN(net243645) );
  NOR2_X2 U5227 ( .A1(n4190), .A2(n4183), .ZN(net243862) );
  AND2_X2 U5228 ( .A1(net243776), .A2(net243775), .ZN(n4190) );
  XNOR2_X2 U5229 ( .A(n4185), .B(net243865), .ZN(net243861) );
  NAND2_X4 U5230 ( .A1(net243780), .A2(net243781), .ZN(net243865) );
  XNOR2_X2 U5231 ( .A(net247850), .B(net243777), .ZN(n4185) );
  INV_X4 U5232 ( .A(net243779), .ZN(net247850) );
  INV_X2 U5233 ( .A(net247850), .ZN(net249128) );
  XNOR2_X2 U5234 ( .A(net243874), .B(net248443), .ZN(net243779) );
  XNOR2_X1 U5235 ( .A(net243875), .B(n4186), .ZN(net248443) );
  XNOR2_X2 U5236 ( .A(net243875), .B(n4186), .ZN(net248442) );
  OAI21_X4 U5237 ( .B1(n4188), .B2(n4187), .A(n4189), .ZN(net243789) );
  INV_X4 U5238 ( .A(net244008), .ZN(n4189) );
  XNOR2_X2 U5239 ( .A(n4189), .B(net244056), .ZN(net244055) );
  INV_X4 U5240 ( .A(net244006), .ZN(n4187) );
  INV_X4 U5241 ( .A(net244005), .ZN(n4188) );
  NAND2_X2 U5242 ( .A1(b[15]), .A2(net246772), .ZN(net243790) );
  NAND2_X4 U5243 ( .A1(net242072), .A2(net242071), .ZN(net241608) );
  INV_X4 U5244 ( .A(net241613), .ZN(net242071) );
  XNOR2_X2 U5245 ( .A(net242072), .B(net242322), .ZN(net242151) );
  NAND2_X4 U5246 ( .A1(net246544), .A2(net246543), .ZN(net246560) );
  NAND2_X4 U5247 ( .A1(net246568), .A2(net246538), .ZN(net246544) );
  INV_X4 U5248 ( .A(net246544), .ZN(net246542) );
  XNOR2_X2 U5249 ( .A(net249149), .B(net246541), .ZN(net246568) );
  NAND2_X4 U5250 ( .A1(n4191), .A2(net246561), .ZN(net246543) );
  NOR2_X1 U5251 ( .A1(net246566), .A2(net245422), .ZN(net246561) );
  INV_X4 U5252 ( .A(n4192), .ZN(n4191) );
  MUX2_X2 U5253 ( .A(net245524), .B(net245525), .S(n4033), .Z(net245523) );
  XNOR2_X2 U5254 ( .A(n4193), .B(net246564), .ZN(n4192) );
  NAND3_X4 U5255 ( .A1(a[30]), .A2(n4194), .A3(b[30]), .ZN(n4193) );
  NAND2_X4 U5256 ( .A1(b[31]), .A2(a[31]), .ZN(n4194) );
  INV_X2 U5257 ( .A(net249149), .ZN(net247741) );
  INV_X4 U5258 ( .A(net246541), .ZN(net246506) );
  OAI22_X1 U5259 ( .A1(n4022), .A2(net246958), .B1(net246770), .B2(net245318), 
        .ZN(net245348) );
  NAND2_X2 U5260 ( .A1(net246539), .A2(n4022), .ZN(net246538) );
  INV_X4 U5261 ( .A(net246566), .ZN(net246577) );
  OAI21_X2 U5262 ( .B1(net246916), .B2(net246579), .A(net246564), .ZN(
        net246578) );
  NAND3_X4 U5263 ( .A1(n4195), .A2(n4197), .A3(n4196), .ZN(net243994) );
  NAND2_X2 U5264 ( .A1(n3967), .A2(net244161), .ZN(n4196) );
  NAND2_X2 U5265 ( .A1(n3967), .A2(net244160), .ZN(n4195) );
  XNOR2_X2 U5266 ( .A(net244160), .B(n3967), .ZN(net244263) );
  INV_X4 U5267 ( .A(net246770), .ZN(net246766) );
  NAND2_X2 U5268 ( .A1(net244160), .A2(net244161), .ZN(n4197) );
  INV_X4 U5269 ( .A(net244163), .ZN(net244160) );
  XNOR2_X2 U5270 ( .A(net244269), .B(net244151), .ZN(net244163) );
  OAI22_X4 U5271 ( .A1(net244378), .A2(net244379), .B1(net247924), .B2(
        net244153), .ZN(net244269) );
  NAND2_X1 U5272 ( .A1(net244153), .A2(net247924), .ZN(net244152) );
  NOR2_X2 U5273 ( .A1(net244154), .A2(net244153), .ZN(net244150) );
  INV_X4 U5274 ( .A(net244154), .ZN(net244378) );
  NAND2_X4 U5275 ( .A1(n4200), .A2(n4201), .ZN(net244161) );
  XNOR2_X2 U5276 ( .A(net244263), .B(net244161), .ZN(net244173) );
  NAND2_X2 U5277 ( .A1(n4199), .A2(net244258), .ZN(n4201) );
  INV_X4 U5278 ( .A(net244260), .ZN(n4199) );
  AOI22_X1 U5279 ( .A1(n4198), .A2(net244260), .B1(n4199), .B2(net244262), 
        .ZN(net244256) );
  AOI21_X4 U5280 ( .B1(net249187), .B2(net244262), .A(n4202), .ZN(n4200) );
  NOR2_X4 U5281 ( .A1(n4198), .A2(net244260), .ZN(n4202) );
  INV_X8 U5282 ( .A(net244262), .ZN(n4198) );
  NAND2_X4 U5283 ( .A1(b[31]), .A2(a[26]), .ZN(net249177) );
  XNOR2_X2 U5284 ( .A(net244270), .B(net248551), .ZN(net244151) );
  INV_X4 U5285 ( .A(net246000), .ZN(net245901) );
  XNOR2_X2 U5286 ( .A(net246109), .B(net246108), .ZN(net246198) );
  AND3_X4 U5287 ( .A1(net246000), .A2(net246002), .A3(net249274), .ZN(
        net248132) );
  NAND2_X4 U5288 ( .A1(b[30]), .A2(a[27]), .ZN(net245250) );
  NAND2_X2 U5289 ( .A1(net242323), .A2(net242324), .ZN(net241612) );
  INV_X4 U5290 ( .A(net242367), .ZN(net242323) );
  NAND2_X2 U5291 ( .A1(net242324), .A2(net242323), .ZN(net242102) );
  XNOR2_X2 U5292 ( .A(net243782), .B(net243401), .ZN(net243651) );
  XNOR2_X2 U5293 ( .A(net243782), .B(net243401), .ZN(net248477) );
  NAND2_X1 U5294 ( .A1(n4203), .A2(net243784), .ZN(net243408) );
  INV_X4 U5295 ( .A(net243785), .ZN(n4203) );
  INV_X4 U5296 ( .A(net243790), .ZN(net243999) );
  INV_X2 U5297 ( .A(net243791), .ZN(net243996) );
  INV_X4 U5298 ( .A(net243784), .ZN(net243998) );
  NAND2_X4 U5299 ( .A1(net245744), .A2(n4204), .ZN(net245691) );
  NAND2_X4 U5300 ( .A1(net245691), .A2(net248865), .ZN(net245680) );
  INV_X4 U5301 ( .A(net245686), .ZN(net245751) );
  NAND3_X2 U5302 ( .A1(net245689), .A2(net249331), .A3(net245751), .ZN(
        net248865) );
  NAND3_X2 U5303 ( .A1(net245689), .A2(net249331), .A3(net245751), .ZN(
        net245742) );
  NOR2_X2 U5304 ( .A1(net248207), .A2(net248867), .ZN(n4205) );
  NAND2_X1 U5305 ( .A1(net248207), .A2(net245750), .ZN(net245960) );
  INV_X1 U5306 ( .A(n4207), .ZN(net248867) );
  INV_X4 U5307 ( .A(net245750), .ZN(n4207) );
  NAND2_X4 U5308 ( .A1(net245962), .A2(n4207), .ZN(net245690) );
  INV_X4 U5309 ( .A(net245745), .ZN(net245744) );
  XNOR2_X2 U5310 ( .A(net245890), .B(net248612), .ZN(net245745) );
  CLKBUF_X3 U5311 ( .A(net245756), .Z(net248612) );
  XNOR2_X2 U5312 ( .A(net245757), .B(net245759), .ZN(net245890) );
  OAI21_X4 U5313 ( .B1(net245985), .B2(n4208), .A(n4212), .ZN(net245750) );
  XNOR2_X2 U5314 ( .A(net245750), .B(net248207), .ZN(net245984) );
  INV_X4 U5315 ( .A(n4211), .ZN(n4212) );
  INV_X8 U5316 ( .A(n4209), .ZN(n4211) );
  AOI21_X4 U5317 ( .B1(n4210), .B2(net247630), .A(n4211), .ZN(net246096) );
  OAI21_X4 U5318 ( .B1(net245989), .B2(net245988), .A(n3957), .ZN(n4209) );
  NOR3_X2 U5319 ( .A1(net245989), .A2(net245988), .A3(n3957), .ZN(n4208) );
  NOR2_X2 U5320 ( .A1(n3957), .A2(net245989), .ZN(n4210) );
  AOI21_X4 U5321 ( .B1(net246581), .B2(net246582), .A(net246910), .ZN(
        net249149) );
  INV_X8 U5322 ( .A(b[30]), .ZN(net246910) );
  AOI21_X2 U5323 ( .B1(net246581), .B2(n4086), .A(net246910), .ZN(net246540)
         );
  NAND2_X4 U5324 ( .A1(a[28]), .A2(b[31]), .ZN(net246541) );
  XNOR2_X2 U5325 ( .A(net246576), .B(net246539), .ZN(net246552) );
  OAI21_X4 U5326 ( .B1(n4213), .B2(n4214), .A(n4215), .ZN(net243313) );
  NAND2_X1 U5327 ( .A1(n4216), .A2(net243367), .ZN(n4215) );
  INV_X4 U5328 ( .A(net243368), .ZN(n4216) );
  NOR2_X2 U5329 ( .A1(n4216), .A2(net243367), .ZN(n4214) );
  XNOR2_X2 U5330 ( .A(net243631), .B(net243630), .ZN(n4213) );
  INV_X4 U5331 ( .A(net243371), .ZN(net243631) );
  XNOR2_X2 U5332 ( .A(net243631), .B(net243630), .ZN(net248988) );
  NAND2_X4 U5333 ( .A1(net247918), .A2(net247919), .ZN(net242832) );
  NAND2_X2 U5334 ( .A1(net247916), .A2(net247917), .ZN(net247919) );
  INV_X1 U5335 ( .A(net242828), .ZN(net247917) );
  INV_X2 U5336 ( .A(net242901), .ZN(net247916) );
  NAND2_X1 U5337 ( .A1(net242901), .A2(net242828), .ZN(net247918) );
  XNOR2_X2 U5338 ( .A(n4218), .B(net242811), .ZN(net242828) );
  NAND2_X2 U5339 ( .A1(net242827), .A2(net242828), .ZN(net242594) );
  OAI21_X4 U5340 ( .B1(net242822), .B2(n4217), .A(net242823), .ZN(n4220) );
  INV_X8 U5341 ( .A(n4221), .ZN(n4217) );
  OAI21_X4 U5342 ( .B1(n4217), .B2(net242817), .A(net242818), .ZN(net242812)
         );
  NAND2_X4 U5343 ( .A1(net243104), .A2(net243105), .ZN(n4221) );
  INV_X4 U5344 ( .A(net243119), .ZN(net243105) );
  NAND3_X2 U5345 ( .A1(net248987), .A2(net243179), .A3(net243105), .ZN(
        net243118) );
  INV_X2 U5346 ( .A(net243106), .ZN(net243104) );
  INV_X4 U5347 ( .A(net248400), .ZN(net242822) );
  XNOR2_X2 U5348 ( .A(net242822), .B(net243177), .ZN(net243176) );
  NAND2_X2 U5349 ( .A1(net242822), .A2(net242823), .ZN(net242819) );
  XNOR2_X2 U5350 ( .A(net243187), .B(n4219), .ZN(net248400) );
  AOI22_X4 U5351 ( .A1(n4039), .A2(net242825), .B1(net242829), .B2(net242830), 
        .ZN(net242901) );
  INV_X8 U5352 ( .A(net242826), .ZN(net242829) );
  NAND2_X2 U5353 ( .A1(net242830), .A2(net242829), .ZN(net242827) );
  INV_X4 U5354 ( .A(net242830), .ZN(net242825) );
  NAND2_X4 U5355 ( .A1(net245952), .A2(net245953), .ZN(net245757) );
  OAI21_X4 U5356 ( .B1(net245955), .B2(net245954), .A(net245956), .ZN(
        net245952) );
  XNOR2_X1 U5357 ( .A(net245773), .B(net245993), .ZN(net245992) );
  INV_X4 U5358 ( .A(net246082), .ZN(net245954) );
  NAND2_X4 U5359 ( .A1(net245955), .A2(net245954), .ZN(net245953) );
  NAND2_X4 U5360 ( .A1(net245953), .A2(net246080), .ZN(net245991) );
  NAND3_X4 U5361 ( .A1(n4224), .A2(n4226), .A3(n4225), .ZN(net245955) );
  NAND2_X2 U5362 ( .A1(n4228), .A2(net249335), .ZN(n4225) );
  INV_X4 U5363 ( .A(net246089), .ZN(n4228) );
  INV_X8 U5364 ( .A(net246105), .ZN(n4229) );
  OAI21_X4 U5365 ( .B1(n4229), .B2(net249076), .A(net246100), .ZN(net249335)
         );
  NAND2_X4 U5366 ( .A1(net247804), .A2(n4229), .ZN(net247807) );
  XNOR2_X2 U5367 ( .A(net246005), .B(n4222), .ZN(net248357) );
  INV_X4 U5368 ( .A(n4223), .ZN(n4222) );
  OAI21_X4 U5369 ( .B1(n4222), .B2(net245907), .A(net245909), .ZN(net245786)
         );
  XNOR2_X2 U5370 ( .A(net246006), .B(net245802), .ZN(n4223) );
  NAND2_X2 U5371 ( .A1(b[5]), .A2(net246772), .ZN(net241003) );
  OAI21_X4 U5372 ( .B1(net241005), .B2(net241006), .A(net241007), .ZN(
        net241002) );
  XOR2_X2 U5373 ( .A(net241006), .B(net241039), .Z(net249059) );
  NAND2_X2 U5374 ( .A1(net246004), .A2(net248623), .ZN(net246000) );
  NAND2_X2 U5375 ( .A1(a[28]), .A2(b[24]), .ZN(net246111) );
  OAI21_X4 U5376 ( .B1(net246199), .B2(net246200), .A(net246201), .ZN(
        net246109) );
  NOR2_X2 U5377 ( .A1(net248925), .A2(n4230), .ZN(net246200) );
  NAND2_X2 U5378 ( .A1(net246204), .A2(net246205), .ZN(n4230) );
  XNOR2_X2 U5379 ( .A(net246199), .B(net246258), .ZN(net246190) );
  NAND2_X2 U5380 ( .A1(net246201), .A2(n4231), .ZN(net246258) );
  OAI21_X4 U5381 ( .B1(net246261), .B2(net248925), .A(net246262), .ZN(
        net246201) );
  NAND3_X4 U5382 ( .A1(net246205), .A2(net246204), .A3(net246260), .ZN(n4231)
         );
  INV_X4 U5383 ( .A(net246204), .ZN(net246262) );
  INV_X4 U5384 ( .A(net246205), .ZN(net246261) );
  INV_X8 U5385 ( .A(net244694), .ZN(net244698) );
  NAND2_X4 U5386 ( .A1(net245678), .A2(net245679), .ZN(net245677) );
  INV_X4 U5387 ( .A(net245680), .ZN(net245678) );
  XNOR2_X2 U5388 ( .A(net245680), .B(net245679), .ZN(net245741) );
  NAND3_X2 U5389 ( .A1(n4232), .A2(net245960), .A3(net245686), .ZN(net245959)
         );
  NAND2_X2 U5390 ( .A1(net248639), .A2(net245690), .ZN(n4232) );
  OAI21_X4 U5391 ( .B1(net244372), .B2(net244373), .A(net244374), .ZN(
        net244136) );
  XNOR2_X2 U5392 ( .A(n4233), .B(n4235), .ZN(net244289) );
  CLKBUF_X3 U5393 ( .A(net244368), .Z(n4235) );
  XNOR2_X2 U5394 ( .A(n4234), .B(net244371), .ZN(n4233) );
  INV_X8 U5395 ( .A(net244369), .ZN(n4234) );
  NAND2_X2 U5396 ( .A1(net246836), .A2(a[24]), .ZN(net244146) );
  NOR2_X4 U5397 ( .A1(net244285), .A2(net244146), .ZN(net244278) );
  INV_X32 U5398 ( .A(a[24]), .ZN(net246756) );
  OAI22_X4 U5399 ( .A1(net246007), .A2(net246008), .B1(n4236), .B2(net246756), 
        .ZN(net246006) );
  INV_X4 U5400 ( .A(net245918), .ZN(n4236) );
  NAND2_X4 U5401 ( .A1(b[22]), .A2(net246772), .ZN(net245686) );
  NAND2_X4 U5402 ( .A1(net249300), .A2(net245960), .ZN(net245689) );
  OAI21_X4 U5403 ( .B1(n4237), .B2(net246386), .A(net246385), .ZN(net246437)
         );
  INV_X1 U5404 ( .A(net246384), .ZN(n4237) );
  XNOR2_X2 U5405 ( .A(n4240), .B(n4241), .ZN(net246396) );
  AOI21_X4 U5406 ( .B1(net246432), .B2(n4243), .A(n4242), .ZN(n4241) );
  INV_X4 U5407 ( .A(net246345), .ZN(n4242) );
  INV_X1 U5408 ( .A(n4239), .ZN(n4243) );
  OAI21_X4 U5409 ( .B1(net246431), .B2(n4239), .A(net246345), .ZN(net246349)
         );
  XNOR2_X2 U5410 ( .A(n4238), .B(net246342), .ZN(n4240) );
  INV_X4 U5411 ( .A(net246346), .ZN(n4238) );
  NAND2_X4 U5412 ( .A1(n4238), .A2(net246349), .ZN(net246353) );
  NAND2_X2 U5413 ( .A1(b[27]), .A2(a[28]), .ZN(net246400) );
  XNOR2_X2 U5414 ( .A(net246206), .B(n4244), .ZN(net248623) );
  INV_X4 U5415 ( .A(net249302), .ZN(n4244) );
  OAI21_X2 U5416 ( .B1(n4244), .B2(net246114), .A(net246071), .ZN(net246113)
         );
  XNOR2_X2 U5417 ( .A(net246206), .B(n4244), .ZN(net246003) );
  AOI22_X4 U5418 ( .A1(n4245), .A2(net246116), .B1(n4253), .B2(net246120), 
        .ZN(net246206) );
  INV_X4 U5419 ( .A(net246116), .ZN(n4253) );
  INV_X4 U5420 ( .A(net246120), .ZN(n4245) );
  NAND2_X2 U5421 ( .A1(n4245), .A2(net246116), .ZN(net246071) );
  XNOR2_X2 U5422 ( .A(n4249), .B(n4248), .ZN(net249302) );
  NAND2_X2 U5423 ( .A1(net249302), .A2(net246077), .ZN(net246070) );
  INV_X4 U5424 ( .A(n4254), .ZN(n4248) );
  NAND2_X4 U5425 ( .A1(net246179), .A2(n4248), .ZN(net246016) );
  XNOR2_X2 U5426 ( .A(n4250), .B(n4255), .ZN(n4254) );
  XOR2_X1 U5427 ( .A(net246132), .B(net246172), .Z(n4255) );
  AOI22_X2 U5428 ( .A1(n4251), .A2(net246127), .B1(n4246), .B2(net246135), 
        .ZN(n4250) );
  INV_X4 U5429 ( .A(net246127), .ZN(n4246) );
  NAND2_X4 U5430 ( .A1(n4246), .A2(net246135), .ZN(net246034) );
  INV_X2 U5431 ( .A(net246135), .ZN(n4251) );
  XNOR2_X2 U5432 ( .A(n4252), .B(n4247), .ZN(n4249) );
  INV_X4 U5433 ( .A(net245429), .ZN(n4247) );
  NAND2_X2 U5434 ( .A1(net246177), .A2(net246176), .ZN(n4252) );
  XNOR2_X2 U5435 ( .A(n4256), .B(net246113), .ZN(net246002) );
  INV_X2 U5436 ( .A(net246077), .ZN(net246114) );
  XNOR2_X2 U5437 ( .A(net246073), .B(net246074), .ZN(n4256) );
  OAI21_X4 U5438 ( .B1(net240918), .B2(n4259), .A(n4260), .ZN(net240763) );
  NAND3_X1 U5439 ( .A1(net240761), .A2(net240763), .A3(net240762), .ZN(out[0])
         );
  INV_X4 U5440 ( .A(net240763), .ZN(net240774) );
  INV_X4 U5441 ( .A(b[0]), .ZN(n4262) );
  NAND2_X2 U5442 ( .A1(a[0]), .A2(n4262), .ZN(net244873) );
  INV_X32 U5443 ( .A(net246974), .ZN(net246970) );
  INV_X4 U5444 ( .A(n4259), .ZN(n4261) );
  INV_X4 U5445 ( .A(net240916), .ZN(net240918) );
  NAND2_X2 U5446 ( .A1(n4263), .A2(net247048), .ZN(n4259) );
  INV_X16 U5447 ( .A(n4267), .ZN(net247048) );
  INV_X8 U5448 ( .A(n4258), .ZN(n4267) );
  INV_X16 U5449 ( .A(n4267), .ZN(net247049) );
  NAND2_X4 U5450 ( .A1(n4257), .A2(net246932), .ZN(n4258) );
  INV_X32 U5451 ( .A(ALUCtrl[0]), .ZN(net246932) );
  INV_X4 U5452 ( .A(n4265), .ZN(n4257) );
  OAI21_X1 U5453 ( .B1(a[30]), .B2(net246904), .A(n4257), .ZN(n3662) );
  OAI21_X2 U5454 ( .B1(net244874), .B2(net244875), .A(n4257), .ZN(net244862)
         );
  NAND2_X2 U5455 ( .A1(n4264), .A2(net245052), .ZN(n4265) );
  INV_X4 U5456 ( .A(ALUCtrl[2]), .ZN(net245052) );
  INV_X4 U5457 ( .A(n4266), .ZN(n4264) );
  NAND3_X4 U5458 ( .A1(n4264), .A2(a[31]), .A3(net246932), .ZN(net240784) );
  NAND2_X2 U5459 ( .A1(ALUCtrl[2]), .A2(n4264), .ZN(net244867) );
  NAND2_X2 U5460 ( .A1(ALUCtrl[3]), .A2(net244841), .ZN(n4266) );
  INV_X4 U5461 ( .A(ALUCtrl[1]), .ZN(net244841) );
  NAND2_X2 U5462 ( .A1(net240782), .A2(a[0]), .ZN(n4263) );
  XNOR2_X2 U5463 ( .A(net244067), .B(net243988), .ZN(net243995) );
  INV_X4 U5464 ( .A(net243991), .ZN(net243988) );
  NAND2_X4 U5465 ( .A1(net243988), .A2(net247223), .ZN(net249194) );
  NAND2_X2 U5466 ( .A1(net243988), .A2(net247223), .ZN(net243729) );
  XNOR2_X2 U5467 ( .A(net243990), .B(net243734), .ZN(net244067) );
  INV_X4 U5468 ( .A(net243989), .ZN(net243990) );
  XNOR2_X2 U5469 ( .A(net240944), .B(n4269), .ZN(n4268) );
  NOR2_X4 U5470 ( .A1(n4270), .A2(n4271), .ZN(n4269) );
  OAI21_X4 U5471 ( .B1(net240944), .B2(n4270), .A(net240933), .ZN(net240949)
         );
  NAND2_X2 U5472 ( .A1(net240933), .A2(net240934), .ZN(net240932) );
  INV_X4 U5473 ( .A(net240952), .ZN(n4272) );
  NAND2_X4 U5474 ( .A1(n4274), .A2(net240952), .ZN(net240934) );
  INV_X4 U5475 ( .A(net240951), .ZN(n4274) );
  XNOR2_X2 U5476 ( .A(n4104), .B(n4024), .ZN(net240931) );
  XNOR2_X2 U5477 ( .A(n4273), .B(net240956), .ZN(net240954) );
  AOI21_X4 U5478 ( .B1(n4277), .B2(n4032), .A(n4054), .ZN(n4273) );
  XOR2_X2 U5479 ( .A(net241573), .B(n4275), .Z(n4277) );
  INV_X2 U5480 ( .A(n4276), .ZN(n4275) );
  XNOR2_X2 U5481 ( .A(net241573), .B(n4275), .ZN(net240961) );
  AOI21_X4 U5482 ( .B1(net241579), .B2(net242103), .A(n3888), .ZN(net241817)
         );
  INV_X4 U5483 ( .A(net240966), .ZN(net240962) );
  XNOR2_X2 U5484 ( .A(net241023), .B(net241024), .ZN(net240966) );
  INV_X4 U5485 ( .A(net240956), .ZN(net240978) );
  OAI21_X2 U5486 ( .B1(n4007), .B2(net244150), .A(net244152), .ZN(net243989)
         );
  CLKBUF_X3 U5487 ( .A(net244075), .Z(net248551) );
  XNOR2_X2 U5488 ( .A(net244076), .B(net244078), .ZN(net244270) );
  NAND2_X2 U5489 ( .A1(b[24]), .A2(net246768), .ZN(net245897) );
  NAND2_X2 U5490 ( .A1(b[5]), .A2(a[28]), .ZN(net241006) );
  XNOR2_X2 U5491 ( .A(n4279), .B(net241018), .ZN(n4278) );
  INV_X4 U5492 ( .A(net241039), .ZN(net241018) );
  NAND2_X4 U5493 ( .A1(net241022), .A2(net241018), .ZN(net241038) );
  XNOR2_X2 U5494 ( .A(net241022), .B(net241582), .ZN(net241573) );
  INV_X4 U5495 ( .A(net241063), .ZN(net241587) );
  XNOR2_X2 U5496 ( .A(n4029), .B(n4280), .ZN(net241071) );
  INV_X4 U5497 ( .A(net241503), .ZN(n4280) );
  XNOR2_X2 U5498 ( .A(net241628), .B(n4280), .ZN(net248620) );
  OAI21_X4 U5499 ( .B1(net241010), .B2(net241011), .A(n3887), .ZN(net241009)
         );
  INV_X4 U5500 ( .A(net241013), .ZN(net241011) );
  INV_X4 U5501 ( .A(net246523), .ZN(net246452) );
  NAND2_X4 U5502 ( .A1(net246452), .A2(net246450), .ZN(net246447) );
  XNOR2_X2 U5503 ( .A(n4282), .B(n4281), .ZN(net246502) );
  XNOR2_X2 U5504 ( .A(net246446), .B(net245541), .ZN(n4281) );
  CLKBUF_X3 U5505 ( .A(net246445), .Z(n4282) );
  AOI21_X4 U5506 ( .B1(net244558), .B2(net244559), .A(net244560), .ZN(
        net244557) );
  OAI21_X4 U5507 ( .B1(net244555), .B2(n4283), .A(net244557), .ZN(net244553)
         );
  AOI211_X2 U5508 ( .C1(net244562), .C2(net244561), .A(net244564), .B(
        net244563), .ZN(net244560) );
  INV_X4 U5509 ( .A(net244565), .ZN(net244563) );
  INV_X4 U5510 ( .A(net244559), .ZN(net244564) );
  NAND2_X4 U5511 ( .A1(n4284), .A2(net244567), .ZN(net244561) );
  INV_X4 U5512 ( .A(n4285), .ZN(n4284) );
  CLKBUF_X3 U5513 ( .A(n4284), .Z(net247211) );
  NOR2_X4 U5514 ( .A1(n4073), .A2(net244567), .ZN(net244668) );
  INV_X8 U5515 ( .A(n4287), .ZN(n4286) );
  INV_X1 U5516 ( .A(n4286), .ZN(net249328) );
  XNOR2_X2 U5517 ( .A(n4286), .B(net245724), .ZN(net247549) );
  NAND2_X4 U5518 ( .A1(n4286), .A2(net244674), .ZN(net244669) );
  XNOR2_X2 U5519 ( .A(net245730), .B(net245614), .ZN(n4287) );
  INV_X4 U5520 ( .A(net244568), .ZN(net244558) );
  NAND2_X2 U5521 ( .A1(net247164), .A2(net244558), .ZN(n4283) );
  NAND2_X2 U5522 ( .A1(b[20]), .A2(net246768), .ZN(net244559) );
  XNOR2_X2 U5523 ( .A(net244568), .B(net244559), .ZN(net244665) );
  INV_X32 U5524 ( .A(b[20]), .ZN(net246832) );
  INV_X4 U5525 ( .A(net244562), .ZN(net244671) );
  XNOR2_X2 U5526 ( .A(net248389), .B(net245613), .ZN(net245612) );
  NAND2_X1 U5527 ( .A1(net244692), .A2(net244685), .ZN(net245613) );
  NAND2_X4 U5528 ( .A1(net241072), .A2(net241073), .ZN(net241070) );
  XNOR2_X2 U5529 ( .A(net241070), .B(net248620), .ZN(net241069) );
  NAND2_X2 U5530 ( .A1(net246766), .A2(b[7]), .ZN(net241063) );
  NOR2_X4 U5531 ( .A1(n4290), .A2(n4291), .ZN(net243780) );
  NAND2_X2 U5532 ( .A1(net243780), .A2(n4043), .ZN(net243778) );
  NOR2_X4 U5533 ( .A1(n4009), .A2(n4293), .ZN(n4291) );
  OR2_X2 U5534 ( .A1(n4289), .A2(net243761), .ZN(n4293) );
  INV_X4 U5535 ( .A(net243763), .ZN(n4289) );
  NAND2_X4 U5536 ( .A1(n4289), .A2(net243765), .ZN(net243868) );
  NOR2_X4 U5537 ( .A1(net243765), .A2(n4289), .ZN(net248371) );
  INV_X8 U5538 ( .A(n4288), .ZN(net243765) );
  NAND2_X1 U5539 ( .A1(net246760), .A2(net243755), .ZN(n4292) );
  XNOR2_X2 U5540 ( .A(net240936), .B(net240937), .ZN(net240924) );
  XNOR2_X2 U5541 ( .A(net240924), .B(net240925), .ZN(net240916) );
  XNOR2_X2 U5542 ( .A(n4294), .B(net240949), .ZN(net240936) );
  XNOR2_X2 U5543 ( .A(net240975), .B(n4295), .ZN(n4294) );
  XNOR2_X2 U5544 ( .A(n4296), .B(net240999), .ZN(n4295) );
  XNOR2_X1 U5545 ( .A(net241023), .B(net241024), .ZN(net248695) );
  XNOR2_X2 U5546 ( .A(net241026), .B(n4297), .ZN(n4296) );
  OAI21_X2 U5547 ( .B1(net249278), .B2(net241029), .A(net249044), .ZN(n4297)
         );
  INV_X4 U5548 ( .A(net249043), .ZN(net249044) );
  NAND2_X2 U5549 ( .A1(net240992), .A2(net249044), .ZN(net240990) );
  XNOR2_X2 U5550 ( .A(net241033), .B(n4298), .ZN(net241029) );
  INV_X4 U5551 ( .A(n4300), .ZN(n4298) );
  XNOR2_X2 U5552 ( .A(n4298), .B(net240994), .ZN(net240989) );
  XNOR2_X2 U5553 ( .A(net241053), .B(net241052), .ZN(n4300) );
  INV_X4 U5554 ( .A(net240994), .ZN(net241033) );
  AND2_X2 U5555 ( .A1(n4299), .A2(net241032), .ZN(net249278) );
  NAND2_X4 U5556 ( .A1(n4299), .A2(net241032), .ZN(net240992) );
  XNOR2_X2 U5557 ( .A(net246277), .B(net248217), .ZN(net246275) );
  XNOR2_X2 U5558 ( .A(net246275), .B(n3934), .ZN(net246269) );
  INV_X4 U5559 ( .A(net248216), .ZN(net248217) );
  INV_X4 U5560 ( .A(net248217), .ZN(net248350) );
  INV_X4 U5561 ( .A(net246243), .ZN(net248216) );
  XNOR2_X2 U5562 ( .A(n4304), .B(net246281), .ZN(net246248) );
  OAI21_X1 U5563 ( .B1(n4301), .B2(net245459), .A(net246236), .ZN(net246281)
         );
  INV_X4 U5564 ( .A(net246238), .ZN(n4301) );
  XNOR2_X2 U5565 ( .A(net246394), .B(n4301), .ZN(net246359) );
  XNOR2_X2 U5566 ( .A(net246129), .B(net246239), .ZN(n4304) );
  NAND2_X2 U5567 ( .A1(b[27]), .A2(net246772), .ZN(net245459) );
  OAI21_X4 U5568 ( .B1(n4302), .B2(n4303), .A(n4305), .ZN(net246236) );
  NAND2_X2 U5569 ( .A1(net246235), .A2(net246236), .ZN(net246131) );
  NAND2_X2 U5570 ( .A1(net246287), .A2(net246288), .ZN(n4303) );
  NAND2_X2 U5571 ( .A1(net246289), .A2(net245459), .ZN(n4302) );
  XNOR2_X2 U5572 ( .A(net246269), .B(net248923), .ZN(net246199) );
  NOR2_X4 U5573 ( .A1(net247632), .A2(net246862), .ZN(net246381) );
  INV_X32 U5574 ( .A(b[23]), .ZN(net246850) );
  NAND2_X4 U5575 ( .A1(net246081), .A2(net246082), .ZN(net246080) );
  NAND2_X4 U5576 ( .A1(b[18]), .A2(a[24]), .ZN(net243578) );
  XNOR2_X2 U5577 ( .A(net240997), .B(net240994), .ZN(net241023) );
  NAND2_X4 U5578 ( .A1(net240991), .A2(net240992), .ZN(net241024) );
  INV_X32 U5579 ( .A(b[26]), .ZN(net246868) );
  OAI22_X4 U5580 ( .A1(n4307), .A2(net243310), .B1(n4045), .B2(n4306), .ZN(
        net243378) );
  INV_X4 U5581 ( .A(net243310), .ZN(n4306) );
  NAND2_X2 U5582 ( .A1(net243307), .A2(net243308), .ZN(net242917) );
  XNOR2_X2 U5583 ( .A(net243285), .B(n4308), .ZN(net243392) );
  NAND2_X2 U5584 ( .A1(net243082), .A2(net243101), .ZN(n4308) );
  INV_X2 U5585 ( .A(net243100), .ZN(net243285) );
  XNOR2_X2 U5586 ( .A(net243285), .B(net243286), .ZN(net243281) );
  XNOR2_X2 U5587 ( .A(net243579), .B(net243301), .ZN(net243391) );
  XNOR2_X2 U5588 ( .A(net243651), .B(net243652), .ZN(net243295) );
  INV_X4 U5589 ( .A(net243082), .ZN(net243078) );
  NAND2_X2 U5590 ( .A1(net243081), .A2(net243082), .ZN(net243098) );
  NAND2_X2 U5591 ( .A1(net243100), .A2(net243101), .ZN(net243099) );
  OAI21_X1 U5592 ( .B1(net243100), .B2(net243279), .A(net243101), .ZN(
        net243278) );
  INV_X4 U5593 ( .A(net243301), .ZN(net243283) );
  INV_X4 U5594 ( .A(net243300), .ZN(net243299) );
  INV_X4 U5595 ( .A(net243580), .ZN(net243298) );
  OAI21_X4 U5596 ( .B1(net248433), .B2(net243296), .A(net243297), .ZN(
        net243284) );
  XNOR2_X2 U5597 ( .A(net248477), .B(net243652), .ZN(net248444) );
  NAND2_X2 U5598 ( .A1(net241020), .A2(n4035), .ZN(net241767) );
  NAND2_X4 U5599 ( .A1(net241045), .A2(net241021), .ZN(net241581) );
  XNOR2_X2 U5600 ( .A(net245616), .B(net247491), .ZN(net248389) );
  INV_X8 U5601 ( .A(net244696), .ZN(net247491) );
  OAI211_X2 U5602 ( .C1(net244543), .C2(net247491), .A(net244545), .B(
        net244540), .ZN(net244535) );
  NAND2_X4 U5603 ( .A1(net245614), .A2(net245615), .ZN(net244692) );
  INV_X8 U5604 ( .A(net244692), .ZN(net244682) );
  OAI21_X4 U5605 ( .B1(net245734), .B2(n4309), .A(n4310), .ZN(net244685) );
  INV_X2 U5606 ( .A(net244685), .ZN(net244681) );
  INV_X4 U5607 ( .A(net244688), .ZN(n4310) );
  NOR2_X2 U5608 ( .A1(n4309), .A2(n4310), .ZN(net245731) );
  INV_X4 U5609 ( .A(n4311), .ZN(n4309) );
  NAND2_X2 U5610 ( .A1(net245737), .A2(net248083), .ZN(n4311) );
  INV_X4 U5611 ( .A(net245732), .ZN(net245734) );
  INV_X4 U5612 ( .A(net244695), .ZN(net244697) );
  NAND2_X4 U5613 ( .A1(net244698), .A2(net244697), .ZN(net244546) );
  NAND2_X4 U5614 ( .A1(n4314), .A2(n4315), .ZN(net244696) );
  NAND2_X4 U5615 ( .A1(net244696), .A2(net244546), .ZN(net244541) );
  NAND2_X4 U5616 ( .A1(n4312), .A2(n4313), .ZN(n4315) );
  INV_X2 U5617 ( .A(net244701), .ZN(n4313) );
  INV_X2 U5618 ( .A(n4313), .ZN(n4316) );
  INV_X4 U5619 ( .A(net245617), .ZN(n4312) );
  NAND2_X2 U5620 ( .A1(net245617), .A2(n4316), .ZN(n4314) );
  NAND2_X2 U5621 ( .A1(b[16]), .A2(net246766), .ZN(net243777) );
  INV_X4 U5622 ( .A(net243777), .ZN(net243770) );
  NOR3_X4 U5623 ( .A1(n4318), .A2(n4319), .A3(n4320), .ZN(net243875) );
  XNOR2_X2 U5624 ( .A(net243875), .B(n3890), .ZN(net248960) );
  NOR2_X4 U5625 ( .A1(n4317), .A2(n4321), .ZN(n4320) );
  NAND2_X2 U5626 ( .A1(net243726), .A2(a[23]), .ZN(n4321) );
  INV_X32 U5627 ( .A(a[23]), .ZN(net246750) );
  INV_X4 U5628 ( .A(net243734), .ZN(net243726) );
  OAI211_X1 U5629 ( .C1(net243726), .C2(net243727), .A(net243728), .B(a[23]), 
        .ZN(net243725) );
  INV_X8 U5630 ( .A(net243728), .ZN(n4317) );
  NAND2_X1 U5631 ( .A1(n4317), .A2(net243733), .ZN(net243731) );
  OAI211_X4 U5632 ( .C1(n4317), .C2(net243734), .A(net243733), .B(net243729), 
        .ZN(n4322) );
  NOR2_X2 U5633 ( .A1(net249194), .A2(net243733), .ZN(n4319) );
  INV_X8 U5634 ( .A(n4322), .ZN(n4318) );
  INV_X2 U5635 ( .A(net243990), .ZN(net247223) );
  NAND2_X2 U5636 ( .A1(net246878), .A2(net246786), .ZN(net246523) );
  INV_X2 U5637 ( .A(net246792), .ZN(net246786) );
  INV_X32 U5638 ( .A(n4323), .ZN(net246878) );
  INV_X16 U5639 ( .A(b[28]), .ZN(n4323) );
  NAND2_X4 U5640 ( .A1(b[27]), .A2(n4323), .ZN(net241542) );
  INV_X16 U5641 ( .A(b[28]), .ZN(net246886) );
  INV_X16 U5642 ( .A(b[28]), .ZN(net246888) );
  NAND2_X4 U5643 ( .A1(n4326), .A2(n4327), .ZN(net242304) );
  CLKBUF_X2 U5644 ( .A(net242304), .Z(net249183) );
  NAND2_X1 U5645 ( .A1(net242304), .A2(net242305), .ZN(net248509) );
  NAND2_X4 U5646 ( .A1(net242304), .A2(net242305), .ZN(net241831) );
  NAND2_X4 U5647 ( .A1(n4325), .A2(n4324), .ZN(n4327) );
  INV_X4 U5648 ( .A(net248776), .ZN(n4324) );
  INV_X4 U5649 ( .A(net242385), .ZN(n4325) );
  NAND2_X2 U5650 ( .A1(net242385), .A2(net248776), .ZN(n4326) );
  NAND2_X4 U5651 ( .A1(b[9]), .A2(net246772), .ZN(net242321) );
  NAND2_X2 U5652 ( .A1(net246766), .A2(b[14]), .ZN(net243301) );
  NAND2_X2 U5653 ( .A1(net243582), .A2(net243584), .ZN(net243300) );
  NAND2_X2 U5654 ( .A1(b[14]), .A2(net246772), .ZN(net243580) );
  INV_X4 U5655 ( .A(net243583), .ZN(n4328) );
  XNOR2_X2 U5656 ( .A(n4341), .B(net243403), .ZN(net243652) );
  NAND2_X2 U5657 ( .A1(net243406), .A2(net243401), .ZN(net243396) );
  INV_X4 U5658 ( .A(net243401), .ZN(net243399) );
  NAND2_X4 U5659 ( .A1(net243298), .A2(net243584), .ZN(net243583) );
  NAND2_X2 U5660 ( .A1(net249197), .A2(net244695), .ZN(net244540) );
  OAI21_X4 U5661 ( .B1(net244701), .B2(net244702), .A(net247168), .ZN(
        net244529) );
  NAND2_X2 U5662 ( .A1(net244701), .A2(net244702), .ZN(net244528) );
  INV_X2 U5663 ( .A(net245775), .ZN(net245896) );
  INV_X4 U5664 ( .A(net245774), .ZN(net245895) );
  NAND2_X2 U5665 ( .A1(n4332), .A2(n4333), .ZN(n4329) );
  NAND2_X2 U5666 ( .A1(n4330), .A2(n4331), .ZN(n4333) );
  INV_X2 U5667 ( .A(net245762), .ZN(n4331) );
  INV_X4 U5668 ( .A(net245906), .ZN(n4330) );
  NAND2_X2 U5669 ( .A1(net245906), .A2(net245762), .ZN(n4332) );
  NAND2_X2 U5670 ( .A1(net244075), .A2(net244076), .ZN(net244074) );
  NAND2_X2 U5671 ( .A1(net244077), .A2(net244076), .ZN(net244072) );
  INV_X4 U5672 ( .A(net244078), .ZN(net244077) );
  NAND2_X4 U5673 ( .A1(a[25]), .A2(b[30]), .ZN(net245317) );
  NAND2_X2 U5674 ( .A1(net243990), .A2(net243991), .ZN(net243728) );
  CLKBUF_X2 U5675 ( .A(net246251), .Z(net248923) );
  XNOR2_X2 U5676 ( .A(n4334), .B(net246237), .ZN(net246394) );
  INV_X4 U5677 ( .A(net245459), .ZN(net246237) );
  NAND2_X2 U5678 ( .A1(net246237), .A2(net246238), .ZN(net246235) );
  NAND3_X2 U5679 ( .A1(net246401), .A2(net246402), .A3(net246403), .ZN(n4334)
         );
  NAND2_X2 U5680 ( .A1(a[28]), .A2(b[26]), .ZN(net246361) );
  NAND2_X2 U5681 ( .A1(b[26]), .A2(net246786), .ZN(net246390) );
  INV_X32 U5682 ( .A(b[31]), .ZN(net246918) );
  NAND2_X2 U5683 ( .A1(n4335), .A2(n4074), .ZN(n4337) );
  NAND2_X2 U5684 ( .A1(net246569), .A2(net246570), .ZN(n4336) );
  NAND2_X2 U5685 ( .A1(net245805), .A2(net245806), .ZN(net246008) );
  NOR2_X2 U5686 ( .A1(n4338), .A2(net245921), .ZN(net246007) );
  XNOR2_X2 U5687 ( .A(n4339), .B(net245369), .ZN(net246005) );
  NAND2_X2 U5688 ( .A1(net245910), .A2(net245911), .ZN(n4339) );
  OAI21_X4 U5689 ( .B1(net245809), .B2(net245802), .A(net245799), .ZN(
        net245808) );
  OAI21_X4 U5690 ( .B1(net243635), .B2(net243583), .A(net243636), .ZN(
        net243634) );
  NOR2_X4 U5691 ( .A1(net246552), .A2(n4340), .ZN(net247173) );
  NAND2_X1 U5692 ( .A1(net246878), .A2(a[31]), .ZN(n4340) );
  INV_X32 U5693 ( .A(a[31]), .ZN(net246812) );
  NAND2_X2 U5694 ( .A1(net246878), .A2(a[30]), .ZN(net246551) );
  XNOR2_X2 U5695 ( .A(n4341), .B(net243403), .ZN(net243395) );
  XNOR2_X2 U5696 ( .A(net249297), .B(n4342), .ZN(net243108) );
  NAND2_X2 U5697 ( .A1(b[11]), .A2(net246772), .ZN(net242830) );
  NAND2_X2 U5698 ( .A1(net242823), .A2(net243118), .ZN(net243177) );
  NAND2_X2 U5699 ( .A1(net243106), .A2(net243119), .ZN(net242823) );
  CLKBUF_X3 U5700 ( .A(net244384), .Z(net247881) );
  INV_X8 U5701 ( .A(net244553), .ZN(net244274) );
  BUF_X8 U5702 ( .A(net244565), .Z(net247164) );
  NAND2_X4 U5703 ( .A1(net244667), .A2(net247164), .ZN(net244666) );
  OAI22_X4 U5704 ( .A1(net244671), .A2(net247211), .B1(net244671), .B2(
        net244567), .ZN(net244555) );
  INV_X4 U5705 ( .A(net244555), .ZN(net244667) );
  XNOR2_X2 U5706 ( .A(net245611), .B(net244671), .ZN(net244659) );
  NAND2_X2 U5707 ( .A1(net240941), .A2(n4345), .ZN(net240929) );
  NAND2_X1 U5708 ( .A1(a[30]), .A2(b[2]), .ZN(n4345) );
  NAND2_X4 U5709 ( .A1(n4344), .A2(a[30]), .ZN(net240930) );
  INV_X4 U5710 ( .A(net240941), .ZN(n4344) );
  XNOR2_X2 U5711 ( .A(net241772), .B(net241773), .ZN(n4346) );
  XNOR2_X2 U5712 ( .A(net241772), .B(net241773), .ZN(net241044) );
  INV_X4 U5713 ( .A(net244554), .ZN(net244273) );
  NAND2_X1 U5714 ( .A1(net244273), .A2(net244274), .ZN(net244272) );
  NOR2_X2 U5715 ( .A1(net242810), .A2(net242811), .ZN(net242580) );
  INV_X4 U5716 ( .A(net242824), .ZN(net242818) );
  INV_X4 U5717 ( .A(net242611), .ZN(net242604) );
  NAND2_X2 U5718 ( .A1(n4350), .A2(net243292), .ZN(net243082) );
  NOR2_X4 U5719 ( .A1(net243290), .A2(net243291), .ZN(n4350) );
  INV_X4 U5720 ( .A(net243396), .ZN(net243290) );
  NOR3_X4 U5721 ( .A1(net243289), .A2(net243290), .A3(net243291), .ZN(
        net243279) );
  NAND3_X2 U5722 ( .A1(net243293), .A2(net243291), .A3(net243294), .ZN(
        net243101) );
  XNOR2_X2 U5723 ( .A(n4351), .B(n4352), .ZN(net243100) );
  XNOR2_X2 U5724 ( .A(net243270), .B(n4353), .ZN(n4352) );
  NAND2_X4 U5725 ( .A1(net243275), .A2(net243404), .ZN(n4353) );
  XNOR2_X1 U5726 ( .A(net243277), .B(n4354), .ZN(n4351) );
  INV_X4 U5727 ( .A(n4349), .ZN(n4354) );
  OAI21_X4 U5728 ( .B1(net243094), .B2(n4354), .A(net243096), .ZN(net243093)
         );
  INV_X8 U5729 ( .A(n4348), .ZN(n4349) );
  XNOR2_X2 U5730 ( .A(net243277), .B(n4349), .ZN(net243271) );
  NAND2_X4 U5731 ( .A1(n4349), .A2(net248780), .ZN(net243066) );
  XNOR2_X2 U5732 ( .A(net243439), .B(net243261), .ZN(n4348) );
  OAI21_X4 U5733 ( .B1(n4356), .B2(net246514), .A(net246515), .ZN(net246468)
         );
  XNOR2_X2 U5734 ( .A(net246510), .B(net246545), .ZN(n4356) );
  INV_X4 U5735 ( .A(net246534), .ZN(net246510) );
  NAND3_X4 U5736 ( .A1(net249225), .A2(net246509), .A3(net246510), .ZN(
        net246332) );
  XNOR2_X2 U5737 ( .A(net246510), .B(net246545), .ZN(net246513) );
  OAI211_X1 U5738 ( .C1(net246788), .C2(a[31]), .A(a[28]), .B(net249231), .ZN(
        n4355) );
  INV_X16 U5739 ( .A(net246918), .ZN(net249231) );
  NAND2_X2 U5740 ( .A1(net240915), .A2(net240916), .ZN(net240762) );
  INV_X4 U5741 ( .A(b[1]), .ZN(n4357) );
  NAND2_X2 U5742 ( .A1(a[1]), .A2(n4357), .ZN(net245029) );
  NAND2_X2 U5743 ( .A1(net240913), .A2(n4357), .ZN(net240910) );
  NAND2_X2 U5744 ( .A1(a[28]), .A2(b[8]), .ZN(net242314) );
  NAND2_X2 U5745 ( .A1(net242316), .A2(net242314), .ZN(net242315) );
  INV_X4 U5746 ( .A(net242314), .ZN(net242313) );
  INV_X4 U5747 ( .A(net243374), .ZN(net243375) );
  OAI22_X4 U5748 ( .A1(net243373), .A2(net243374), .B1(net243375), .B2(
        net243376), .ZN(net243630) );
  NAND2_X4 U5749 ( .A1(net243371), .A2(n4359), .ZN(net243185) );
  NAND2_X2 U5750 ( .A1(net243373), .A2(net243374), .ZN(n4359) );
  NAND2_X2 U5751 ( .A1(net246778), .A2(b[4]), .ZN(net240956) );
  OAI211_X2 U5752 ( .C1(net241563), .C2(n4360), .A(net241565), .B(net241566), 
        .ZN(net240958) );
  OAI21_X2 U5753 ( .B1(net241562), .B2(net240986), .A(net240958), .ZN(
        net241561) );
  INV_X4 U5754 ( .A(net241567), .ZN(n4360) );
  XNOR2_X2 U5755 ( .A(net241767), .B(net249059), .ZN(net241582) );
  XNOR2_X2 U5756 ( .A(n4361), .B(net242074), .ZN(net241607) );
  NAND2_X4 U5757 ( .A1(net241600), .A2(net242076), .ZN(n4361) );
  XNOR2_X2 U5758 ( .A(n4362), .B(net242074), .ZN(net242097) );
  NAND2_X2 U5759 ( .A1(net241600), .A2(net242076), .ZN(n4362) );
  NAND2_X2 U5760 ( .A1(net241599), .A2(net241600), .ZN(net241625) );
  NAND2_X4 U5761 ( .A1(net241599), .A2(net241600), .ZN(net241598) );
  OAI21_X2 U5762 ( .B1(net244687), .B2(net244688), .A(net244684), .ZN(
        net244686) );
  INV_X4 U5763 ( .A(net244684), .ZN(net244683) );
  INV_X32 U5764 ( .A(b[21]), .ZN(net246838) );
  NOR3_X4 U5765 ( .A1(net246091), .A2(net247632), .A3(net246838), .ZN(
        net245981) );
  INV_X32 U5766 ( .A(net246838), .ZN(net246836) );
  AOI21_X4 U5767 ( .B1(n4363), .B2(net242894), .A(n4364), .ZN(net242835) );
  XNOR2_X2 U5768 ( .A(net243175), .B(net243176), .ZN(n4364) );
  INV_X4 U5769 ( .A(net242896), .ZN(n4363) );
  NAND2_X2 U5770 ( .A1(n4365), .A2(net242896), .ZN(net242839) );
  INV_X4 U5771 ( .A(net242894), .ZN(n4365) );
  OAI21_X1 U5772 ( .B1(n4365), .B2(net243166), .A(net242900), .ZN(net243168)
         );
  NOR2_X4 U5773 ( .A1(net243171), .A2(n4365), .ZN(net243172) );
  NOR2_X4 U5774 ( .A1(net242898), .A2(net242894), .ZN(net243164) );
  OAI211_X2 U5775 ( .C1(n4366), .C2(net244177), .A(net244178), .B(n4367), .ZN(
        net243863) );
  NAND2_X2 U5776 ( .A1(net243775), .A2(net243863), .ZN(net244062) );
  INV_X4 U5777 ( .A(net244180), .ZN(n4367) );
  INV_X4 U5778 ( .A(net244181), .ZN(n4366) );
  XNOR2_X2 U5779 ( .A(net244064), .B(net243765), .ZN(net243776) );
  OAI21_X4 U5780 ( .B1(n4368), .B2(n4369), .A(net246272), .ZN(net246251) );
  NAND2_X4 U5781 ( .A1(n3934), .A2(net246251), .ZN(net246118) );
  INV_X2 U5782 ( .A(net246274), .ZN(n4368) );
  NAND2_X4 U5783 ( .A1(net244669), .A2(net244668), .ZN(net244565) );
  NAND2_X2 U5784 ( .A1(net246760), .A2(b[22]), .ZN(net244695) );
  INV_X1 U5785 ( .A(net244287), .ZN(net249352) );
  NAND2_X4 U5786 ( .A1(n8095), .A2(n8097), .ZN(n7814) );
  XNOR2_X2 U5787 ( .A(n4929), .B(n3966), .ZN(n4883) );
  XNOR2_X2 U5788 ( .A(n4370), .B(n7771), .ZN(n8025) );
  XNOR2_X2 U5789 ( .A(n8009), .B(n8010), .ZN(n4370) );
  NAND2_X1 U5790 ( .A1(n8011), .A2(n8012), .ZN(n7771) );
  AND3_X4 U5791 ( .A1(n4877), .A2(n4876), .A3(n4875), .ZN(net249076) );
  NOR2_X2 U5792 ( .A1(n7302), .A2(n4408), .ZN(n7305) );
  INV_X2 U5793 ( .A(n7103), .ZN(n4408) );
  NAND2_X4 U5794 ( .A1(net245739), .A2(net245738), .ZN(net244690) );
  INV_X1 U5795 ( .A(n6651), .ZN(n4371) );
  INV_X2 U5796 ( .A(n4371), .ZN(n4372) );
  AOI22_X2 U5797 ( .A1(net245697), .A2(net245698), .B1(n5087), .B2(net244567), 
        .ZN(net245611) );
  XNOR2_X2 U5798 ( .A(n4471), .B(n8259), .ZN(net241773) );
  INV_X1 U5799 ( .A(net242877), .ZN(net249298) );
  XNOR2_X2 U5800 ( .A(n5123), .B(n5056), .ZN(n4373) );
  INV_X4 U5801 ( .A(n4373), .ZN(n5132) );
  INV_X2 U5802 ( .A(n5121), .ZN(n5123) );
  XNOR2_X2 U5803 ( .A(n4375), .B(n4374), .ZN(n8456) );
  XNOR2_X2 U5804 ( .A(n8446), .B(n8445), .ZN(n4375) );
  OAI21_X2 U5805 ( .B1(n8511), .B2(n8510), .A(n8509), .ZN(n8513) );
  NAND2_X2 U5806 ( .A1(net243395), .A2(net243396), .ZN(net243294) );
  NAND2_X1 U5807 ( .A1(b[6]), .A2(net246766), .ZN(net241032) );
  INV_X4 U5808 ( .A(n4696), .ZN(n4694) );
  AOI22_X4 U5809 ( .A1(n7283), .A2(n7282), .B1(n7287), .B2(n7286), .ZN(n7216)
         );
  INV_X4 U5810 ( .A(n4377), .ZN(n4378) );
  NOR2_X2 U5811 ( .A1(net241757), .A2(net241758), .ZN(n8146) );
  NAND2_X2 U5812 ( .A1(net246407), .A2(n4729), .ZN(net246402) );
  AND2_X2 U5813 ( .A1(n6726), .A2(net243578), .ZN(n4379) );
  NAND2_X4 U5814 ( .A1(net248960), .A2(net249104), .ZN(n6726) );
  INV_X2 U5815 ( .A(n6062), .ZN(n4380) );
  INV_X1 U5816 ( .A(net246071), .ZN(net246075) );
  NAND2_X2 U5817 ( .A1(net249130), .A2(net246525), .ZN(n4495) );
  INV_X2 U5818 ( .A(net248913), .ZN(net246525) );
  NAND2_X4 U5819 ( .A1(n4678), .A2(n5294), .ZN(net249225) );
  INV_X2 U5820 ( .A(n4763), .ZN(n4812) );
  INV_X2 U5821 ( .A(net246792), .ZN(net246790) );
  OAI21_X4 U5822 ( .B1(n5069), .B2(n5070), .A(n5068), .ZN(n5085) );
  XNOR2_X2 U5823 ( .A(net244457), .B(net247881), .ZN(net249187) );
  INV_X8 U5824 ( .A(net249177), .ZN(net247778) );
  INV_X8 U5825 ( .A(b[31]), .ZN(net246920) );
  XNOR2_X2 U5826 ( .A(n4383), .B(n4384), .ZN(n6486) );
  XNOR2_X2 U5827 ( .A(n6477), .B(n6475), .ZN(n4383) );
  OAI21_X4 U5828 ( .B1(net245782), .B2(net245783), .A(n4031), .ZN(n5058) );
  NAND2_X2 U5829 ( .A1(n4730), .A2(n4729), .ZN(net246403) );
  CLKBUF_X3 U5830 ( .A(n6185), .Z(n4385) );
  INV_X2 U5831 ( .A(net242379), .ZN(net242658) );
  XNOR2_X2 U5832 ( .A(n4387), .B(n6795), .ZN(n4386) );
  INV_X4 U5833 ( .A(n4386), .ZN(n6802) );
  XNOR2_X2 U5834 ( .A(n6793), .B(n6792), .ZN(n4387) );
  NOR2_X2 U5835 ( .A1(n8467), .A2(n8466), .ZN(n8470) );
  CLKBUF_X2 U5836 ( .A(n6772), .Z(n4388) );
  XNOR2_X2 U5837 ( .A(n6364), .B(n3968), .ZN(n4470) );
  NAND2_X2 U5838 ( .A1(net243399), .A2(net243400), .ZN(net243293) );
  NOR2_X2 U5839 ( .A1(net244682), .A2(net244686), .ZN(n5933) );
  XNOR2_X2 U5840 ( .A(n4390), .B(n4389), .ZN(n7145) );
  XNOR2_X2 U5841 ( .A(n7135), .B(n7134), .ZN(n4390) );
  INV_X4 U5842 ( .A(net243747), .ZN(net249104) );
  INV_X1 U5843 ( .A(n6332), .ZN(n4391) );
  XNOR2_X2 U5844 ( .A(n4393), .B(n4394), .ZN(n7471) );
  XNOR2_X2 U5845 ( .A(n7477), .B(n7480), .ZN(n4393) );
  NAND2_X4 U5846 ( .A1(n6684), .A2(net248403), .ZN(net243582) );
  NAND2_X2 U5847 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  INV_X1 U5848 ( .A(n4785), .ZN(n4395) );
  XOR2_X2 U5849 ( .A(n5009), .B(n5008), .Z(n4396) );
  INV_X2 U5850 ( .A(net243639), .ZN(net248403) );
  AOI21_X2 U5851 ( .B1(n6730), .B2(n6728), .A(n6727), .ZN(n6732) );
  NAND2_X1 U5852 ( .A1(net243172), .A2(net242899), .ZN(n7021) );
  OAI221_X4 U5853 ( .B1(n4928), .B2(net245921), .C1(n4927), .C2(net245921), 
        .A(n4926), .ZN(net245918) );
  INV_X2 U5854 ( .A(net244173), .ZN(net244244) );
  NOR2_X2 U5855 ( .A1(n5446), .A2(n5445), .ZN(n5465) );
  NAND2_X4 U5856 ( .A1(n6530), .A2(n6529), .ZN(net243763) );
  NOR2_X2 U5857 ( .A1(n6510), .A2(n6509), .ZN(n6513) );
  XNOR2_X2 U5858 ( .A(n4910), .B(n3956), .ZN(n4397) );
  XNOR2_X2 U5859 ( .A(n6870), .B(n6609), .ZN(n4398) );
  INV_X8 U5860 ( .A(n5004), .ZN(n5006) );
  OAI211_X4 U5861 ( .C1(n4841), .C2(n4840), .A(n4839), .B(net246133), .ZN(
        n4885) );
  NAND2_X1 U5862 ( .A1(n3983), .A2(n7622), .ZN(n7625) );
  XNOR2_X2 U5863 ( .A(n8165), .B(n8079), .ZN(n4399) );
  NAND2_X2 U5864 ( .A1(net241563), .A2(net241565), .ZN(net240985) );
  NOR2_X2 U5865 ( .A1(n6439), .A2(n4466), .ZN(n6442) );
  NOR2_X2 U5866 ( .A1(n8478), .A2(n8477), .ZN(n8481) );
  XNOR2_X2 U5867 ( .A(n7698), .B(n7785), .ZN(n4400) );
  NAND2_X4 U5868 ( .A1(n5012), .A2(n5011), .ZN(n5021) );
  AOI21_X2 U5869 ( .B1(net247778), .B2(n4766), .A(net246327), .ZN(n4768) );
  CLKBUF_X3 U5870 ( .A(n5865), .Z(n4401) );
  INV_X2 U5871 ( .A(net249187), .ZN(net244257) );
  XNOR2_X1 U5872 ( .A(n6257), .B(n4378), .ZN(n6388) );
  NAND2_X2 U5873 ( .A1(n6666), .A2(n6665), .ZN(n6747) );
  INV_X4 U5874 ( .A(net248693), .ZN(net242899) );
  NAND2_X1 U5875 ( .A1(net243164), .A2(net248693), .ZN(n7019) );
  INV_X2 U5876 ( .A(n4811), .ZN(n4791) );
  XNOR2_X2 U5877 ( .A(n5139), .B(net248449), .ZN(n4403) );
  INV_X2 U5878 ( .A(net244655), .ZN(net248449) );
  OAI21_X1 U5879 ( .B1(n8725), .B2(n8724), .A(n8723), .ZN(n8726) );
  NAND2_X4 U5880 ( .A1(net248040), .A2(n4477), .ZN(net243175) );
  INV_X2 U5881 ( .A(n7622), .ZN(n7385) );
  NOR2_X2 U5882 ( .A1(n6336), .A2(n6170), .ZN(n6207) );
  NAND2_X2 U5883 ( .A1(n4385), .A2(n6184), .ZN(n6186) );
  NOR2_X2 U5884 ( .A1(n4385), .A2(n6184), .ZN(n6188) );
  XNOR2_X2 U5885 ( .A(n4809), .B(n4792), .ZN(n4404) );
  INV_X1 U5886 ( .A(n4761), .ZN(n4762) );
  INV_X2 U5887 ( .A(n6051), .ZN(n4405) );
  INV_X4 U5888 ( .A(n4405), .ZN(n4406) );
  XNOR2_X2 U5889 ( .A(n8144), .B(n8145), .ZN(n4407) );
  INV_X2 U5890 ( .A(net247821), .ZN(net248893) );
  NAND2_X1 U5891 ( .A1(n7881), .A2(n7880), .ZN(n7883) );
  NAND2_X4 U5892 ( .A1(n7690), .A2(n7689), .ZN(n7880) );
  OAI21_X4 U5893 ( .B1(n4464), .B2(n6385), .A(net244006), .ZN(net244056) );
  NAND2_X4 U5894 ( .A1(n6076), .A2(n6075), .ZN(n6195) );
  INV_X2 U5895 ( .A(n7226), .ZN(n7225) );
  NAND2_X2 U5896 ( .A1(net242916), .A2(net242917), .ZN(n7226) );
  XNOR2_X2 U5897 ( .A(net246445), .B(net248353), .ZN(n4706) );
  INV_X4 U5898 ( .A(n5909), .ZN(n4409) );
  INV_X1 U5899 ( .A(n5046), .ZN(n4410) );
  CLKBUF_X3 U5900 ( .A(n6946), .Z(n4417) );
  XNOR2_X2 U5901 ( .A(n4760), .B(n4840), .ZN(n4411) );
  NAND2_X4 U5902 ( .A1(n4803), .A2(n4804), .ZN(n4760) );
  INV_X2 U5903 ( .A(n4725), .ZN(n4412) );
  INV_X4 U5904 ( .A(n4890), .ZN(n4413) );
  INV_X4 U5905 ( .A(n4413), .ZN(n4414) );
  XNOR2_X2 U5906 ( .A(n5119), .B(n4420), .ZN(n4415) );
  NAND2_X2 U5907 ( .A1(n4942), .A2(n4941), .ZN(n5068) );
  XNOR2_X2 U5908 ( .A(n4085), .B(n4723), .ZN(n4416) );
  NAND2_X2 U5909 ( .A1(net245959), .A2(net245742), .ZN(n4974) );
  NAND2_X2 U5910 ( .A1(n4976), .A2(n4975), .ZN(n4936) );
  NAND2_X4 U5911 ( .A1(n7220), .A2(n7219), .ZN(n7275) );
  AOI21_X4 U5912 ( .B1(a[18]), .B2(net246878), .A(n5869), .ZN(n4439) );
  INV_X2 U5913 ( .A(n5029), .ZN(n4953) );
  OAI22_X4 U5914 ( .A1(n6594), .A2(n6593), .B1(n6592), .B2(n6591), .ZN(n6544)
         );
  NAND2_X4 U5915 ( .A1(n6598), .A2(n6597), .ZN(n6874) );
  XNOR2_X2 U5916 ( .A(n4824), .B(n4825), .ZN(n4440) );
  NAND2_X1 U5917 ( .A1(b[23]), .A2(a[30]), .ZN(n4822) );
  INV_X4 U5918 ( .A(n6667), .ZN(n4418) );
  NAND3_X2 U5919 ( .A1(n6842), .A2(n6841), .A3(n6840), .ZN(n7003) );
  OAI21_X2 U5920 ( .B1(n4435), .B2(n6835), .A(n6834), .ZN(n6840) );
  NOR2_X2 U5921 ( .A1(n7072), .A2(n6941), .ZN(n4419) );
  NAND2_X1 U5922 ( .A1(a[23]), .A2(b[16]), .ZN(n7073) );
  INV_X2 U5923 ( .A(n7073), .ZN(n6941) );
  XNOR2_X2 U5924 ( .A(n7441), .B(n7804), .ZN(net248776) );
  NAND2_X4 U5925 ( .A1(n7880), .A2(n7881), .ZN(n7694) );
  NAND2_X1 U5926 ( .A1(n7443), .A2(n7438), .ZN(n7444) );
  INV_X1 U5927 ( .A(n5967), .ZN(n4421) );
  INV_X8 U5928 ( .A(n8082), .ZN(n7796) );
  XNOR2_X2 U5929 ( .A(n6159), .B(n6158), .ZN(n4422) );
  NAND2_X4 U5930 ( .A1(n6304), .A2(n6305), .ZN(n6158) );
  XNOR2_X2 U5931 ( .A(n7165), .B(n4424), .ZN(n6997) );
  NAND2_X4 U5932 ( .A1(net242594), .A2(net242595), .ZN(n7438) );
  NAND3_X2 U5933 ( .A1(n7804), .A2(n7801), .A3(n7803), .ZN(n7811) );
  NAND3_X2 U5934 ( .A1(n7887), .A2(n7886), .A3(n7885), .ZN(n4425) );
  NAND2_X2 U5935 ( .A1(n6244), .A2(n6245), .ZN(n6313) );
  NOR2_X1 U5936 ( .A1(n6248), .A2(n6313), .ZN(n6249) );
  INV_X1 U5937 ( .A(n6108), .ZN(n4427) );
  INV_X4 U5938 ( .A(n6884), .ZN(n6596) );
  INV_X1 U5939 ( .A(n4962), .ZN(n4909) );
  XNOR2_X1 U5940 ( .A(n8724), .B(n8486), .ZN(n4428) );
  NAND2_X4 U5941 ( .A1(n8723), .A2(n8722), .ZN(n8486) );
  INV_X1 U5942 ( .A(n5095), .ZN(n4429) );
  INV_X2 U5943 ( .A(n4429), .ZN(n4430) );
  INV_X4 U5944 ( .A(n8033), .ZN(n4431) );
  INV_X8 U5945 ( .A(n4431), .ZN(n4432) );
  OAI22_X4 U5946 ( .A1(n7606), .A2(n7604), .B1(n7779), .B2(n7780), .ZN(n7695)
         );
  NAND2_X4 U5947 ( .A1(n7603), .A2(n7288), .ZN(n7780) );
  INV_X4 U5948 ( .A(n7217), .ZN(n7222) );
  NOR2_X2 U5949 ( .A1(n3910), .A2(n7865), .ZN(n7867) );
  NAND2_X4 U5950 ( .A1(n7876), .A2(n7877), .ZN(net241600) );
  XNOR2_X2 U5951 ( .A(n4461), .B(n4460), .ZN(n4433) );
  NOR2_X2 U5952 ( .A1(n7637), .A2(n7636), .ZN(n7640) );
  INV_X2 U5953 ( .A(n8080), .ZN(n8090) );
  OAI21_X2 U5954 ( .B1(n7148), .B2(n7147), .A(n7146), .ZN(n7150) );
  NOR2_X2 U5955 ( .A1(n4404), .A2(n4834), .ZN(n4841) );
  INV_X2 U5956 ( .A(n4838), .ZN(n4793) );
  INV_X2 U5957 ( .A(n6244), .ZN(n6242) );
  NAND2_X2 U5958 ( .A1(n6248), .A2(n6313), .ZN(n6312) );
  INV_X2 U5959 ( .A(n6313), .ZN(n6315) );
  NOR2_X2 U5960 ( .A1(n6587), .A2(n6586), .ZN(n6590) );
  NOR2_X2 U5961 ( .A1(n6300), .A2(n6299), .ZN(n6303) );
  INV_X2 U5962 ( .A(n7692), .ZN(n7686) );
  INV_X2 U5963 ( .A(net249300), .ZN(net248639) );
  OAI21_X2 U5964 ( .B1(n8088), .B2(n8087), .A(n8086), .ZN(n8089) );
  OAI21_X4 U5965 ( .B1(n5910), .B2(n5909), .A(n4488), .ZN(n5911) );
  INV_X8 U5966 ( .A(n5128), .ZN(n5910) );
  INV_X4 U5967 ( .A(n6836), .ZN(n6744) );
  XNOR2_X2 U5968 ( .A(n4438), .B(n5900), .ZN(n4437) );
  INV_X4 U5969 ( .A(n4437), .ZN(n5909) );
  XNOR2_X2 U5970 ( .A(n5897), .B(n5898), .ZN(n4438) );
  NOR2_X1 U5971 ( .A1(n7947), .A2(n7946), .ZN(n7950) );
  NAND2_X1 U5972 ( .A1(n7947), .A2(n7946), .ZN(n7948) );
  OAI21_X2 U5973 ( .B1(n4403), .B2(n4053), .A(n6097), .ZN(n6099) );
  XNOR2_X2 U5974 ( .A(n4440), .B(net246188), .ZN(n5411) );
  NAND2_X2 U5975 ( .A1(n8181), .A2(n8180), .ZN(n8183) );
  INV_X2 U5976 ( .A(net246072), .ZN(net248615) );
  INV_X2 U5977 ( .A(net246073), .ZN(net246072) );
  NAND2_X2 U5978 ( .A1(net247820), .A2(net247821), .ZN(n4500) );
  XNOR2_X2 U5979 ( .A(n4982), .B(n4981), .ZN(n4449) );
  OAI22_X4 U5980 ( .A1(n4998), .A2(n4997), .B1(n4996), .B2(n4995), .ZN(n5009)
         );
  INV_X4 U5981 ( .A(net246190), .ZN(net246188) );
  NAND3_X2 U5982 ( .A1(n7379), .A2(n7378), .A3(n7377), .ZN(n7599) );
  XNOR2_X1 U5983 ( .A(n4411), .B(n4793), .ZN(n4441) );
  CLKBUF_X3 U5984 ( .A(n5340), .Z(n4442) );
  NOR3_X2 U5985 ( .A1(net241824), .A2(net241829), .A3(net241749), .ZN(
        net241828) );
  INV_X1 U5986 ( .A(n7769), .ZN(n4443) );
  INV_X4 U5987 ( .A(n4443), .ZN(n4444) );
  NOR2_X2 U5988 ( .A1(n7505), .A2(n3970), .ZN(n4445) );
  INV_X4 U5989 ( .A(n4445), .ZN(n7728) );
  NAND2_X1 U5990 ( .A1(net245741), .A2(net245740), .ZN(n4507) );
  XNOR2_X2 U5991 ( .A(n4449), .B(n4983), .ZN(net248549) );
  NAND2_X4 U5992 ( .A1(n8328), .A2(n8327), .ZN(n8150) );
  INV_X1 U5993 ( .A(n6210), .ZN(n4446) );
  XNOR2_X2 U5994 ( .A(n7059), .B(n7080), .ZN(n7060) );
  NAND2_X1 U5995 ( .A1(net248371), .A2(net246760), .ZN(n6603) );
  NAND2_X2 U5996 ( .A1(n4470), .A2(n6477), .ZN(n6482) );
  BUF_X32 U5997 ( .A(n6545), .Z(n4447) );
  INV_X1 U5998 ( .A(n7400), .ZN(n4448) );
  NAND2_X2 U5999 ( .A1(net244369), .A2(net244368), .ZN(n6329) );
  NAND2_X4 U6000 ( .A1(b[20]), .A2(a[30]), .ZN(n4983) );
  INV_X1 U6001 ( .A(n6688), .ZN(n4450) );
  INV_X16 U6002 ( .A(net246908), .ZN(net248516) );
  INV_X16 U6003 ( .A(net246908), .ZN(net248517) );
  INV_X16 U6004 ( .A(net246908), .ZN(net246902) );
  OAI21_X2 U6005 ( .B1(n3907), .B2(net242882), .A(net242883), .ZN(n7233) );
  NOR2_X2 U6006 ( .A1(n5143), .A2(n5142), .ZN(n5146) );
  INV_X2 U6007 ( .A(net246407), .ZN(net248511) );
  OAI211_X4 U6008 ( .C1(n7813), .C2(n7812), .A(n3980), .B(n7811), .ZN(n8097)
         );
  INV_X1 U6009 ( .A(n7460), .ZN(n7298) );
  NOR2_X2 U6010 ( .A1(n7299), .A2(n7298), .ZN(n7300) );
  INV_X4 U6011 ( .A(n8028), .ZN(n4451) );
  NOR2_X1 U6012 ( .A1(net242066), .A2(net242067), .ZN(n7683) );
  NOR2_X2 U6013 ( .A1(net248788), .A2(net242319), .ZN(n7679) );
  INV_X2 U6014 ( .A(n6471), .ZN(n6469) );
  INV_X2 U6015 ( .A(n6472), .ZN(n6470) );
  XNOR2_X2 U6016 ( .A(n7309), .B(n7203), .ZN(n4452) );
  AOI21_X2 U6017 ( .B1(n4858), .B2(n4521), .A(n4857), .ZN(n4453) );
  OAI21_X4 U6018 ( .B1(n3906), .B2(n6312), .A(net244173), .ZN(n6530) );
  OAI21_X1 U6019 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(n4454) );
  XNOR2_X2 U6020 ( .A(n7007), .B(n4108), .ZN(n4455) );
  NAND2_X2 U6021 ( .A1(n3933), .A2(n5031), .ZN(n5036) );
  INV_X1 U6022 ( .A(n8256), .ZN(n4456) );
  NAND2_X4 U6023 ( .A1(net243096), .A2(net248780), .ZN(net243277) );
  XNOR2_X2 U6024 ( .A(n6079), .B(n6078), .ZN(n4458) );
  OAI21_X2 U6025 ( .B1(net241276), .B2(net248620), .A(net241072), .ZN(n8553)
         );
  AOI21_X1 U6026 ( .B1(n6596), .B2(n6887), .A(n6595), .ZN(n6686) );
  NAND2_X4 U6027 ( .A1(n5082), .A2(n5939), .ZN(n5080) );
  INV_X1 U6028 ( .A(net248444), .ZN(net248432) );
  INV_X2 U6029 ( .A(net248432), .ZN(net248433) );
  NAND2_X4 U6030 ( .A1(n4404), .A2(n4834), .ZN(n4839) );
  XNOR2_X2 U6031 ( .A(n4461), .B(n4460), .ZN(n7518) );
  XNOR2_X2 U6032 ( .A(n7507), .B(n7508), .ZN(n4461) );
  NAND2_X2 U6033 ( .A1(n6099), .A2(n6100), .ZN(n6240) );
  BUF_X4 U6034 ( .A(n7463), .Z(n4462) );
  NAND3_X2 U6035 ( .A1(n6951), .A2(n6950), .A3(n6952), .ZN(n6947) );
  OAI21_X2 U6036 ( .B1(n6876), .B2(n6732), .A(n6862), .ZN(n6946) );
  INV_X4 U6037 ( .A(n4852), .ZN(n4849) );
  XNOR2_X2 U6038 ( .A(n7594), .B(n7593), .ZN(n4463) );
  NAND2_X1 U6039 ( .A1(n7693), .A2(n7692), .ZN(n7881) );
  XNOR2_X2 U6040 ( .A(n6253), .B(net244243), .ZN(n4464) );
  INV_X1 U6041 ( .A(n7370), .ZN(n4465) );
  XNOR2_X2 U6042 ( .A(net245249), .B(net249177), .ZN(net248379) );
  OAI21_X4 U6043 ( .B1(n4791), .B2(n4810), .A(n4808), .ZN(n4792) );
  OAI21_X4 U6044 ( .B1(n4441), .B2(net246130), .A(net246131), .ZN(n4867) );
  CLKBUF_X3 U6045 ( .A(n6438), .Z(n4466) );
  INV_X4 U6046 ( .A(n6734), .ZN(n4467) );
  XNOR2_X2 U6047 ( .A(n7464), .B(n7357), .ZN(n4468) );
  XNOR2_X2 U6048 ( .A(n4453), .B(n4902), .ZN(n4890) );
  INV_X4 U6049 ( .A(net248353), .ZN(net248354) );
  XNOR2_X2 U6050 ( .A(n7388), .B(n7387), .ZN(n4469) );
  INV_X1 U6051 ( .A(net240783), .ZN(net240912) );
  OAI21_X2 U6052 ( .B1(n8860), .B2(n8859), .A(b[1]), .ZN(net240767) );
  XNOR2_X2 U6053 ( .A(n8269), .B(net241625), .ZN(n4471) );
  NOR2_X2 U6054 ( .A1(n8488), .A2(n8487), .ZN(n8491) );
  OAI21_X2 U6055 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n8498) );
  AOI21_X2 U6056 ( .B1(n8495), .B2(n8494), .A(n8496), .ZN(n8174) );
  NAND2_X2 U6057 ( .A1(n8168), .A2(n8169), .ZN(n8066) );
  OAI21_X2 U6058 ( .B1(n4771), .B2(n4713), .A(n4395), .ZN(n4776) );
  OAI22_X2 U6059 ( .A1(n6382), .A2(n6381), .B1(n6384), .B2(n6383), .ZN(n6254)
         );
  NAND2_X4 U6060 ( .A1(n5331), .A2(net246381), .ZN(n4733) );
  INV_X8 U6061 ( .A(n4879), .ZN(n4832) );
  NOR2_X1 U6062 ( .A1(n4012), .A2(n7174), .ZN(n7178) );
  NAND2_X1 U6063 ( .A1(n4012), .A2(n7174), .ZN(n7176) );
  INV_X4 U6064 ( .A(n7823), .ZN(n8104) );
  OAI21_X2 U6065 ( .B1(n4856), .B2(n4855), .A(n4854), .ZN(n4472) );
  NAND2_X1 U6066 ( .A1(n4785), .A2(n4784), .ZN(n4787) );
  INV_X1 U6067 ( .A(net246353), .ZN(net246407) );
  NAND2_X2 U6068 ( .A1(n5062), .A2(n5061), .ZN(n5131) );
  XNOR2_X1 U6069 ( .A(n6733), .B(n6754), .ZN(n6735) );
  NOR2_X4 U6070 ( .A1(n4718), .A2(n4766), .ZN(n4719) );
  INV_X4 U6071 ( .A(n4823), .ZN(n4824) );
  XNOR2_X2 U6072 ( .A(n6746), .B(n6668), .ZN(n6527) );
  NAND2_X2 U6073 ( .A1(n6536), .A2(n6535), .ZN(n6679) );
  NAND2_X1 U6074 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  NAND2_X1 U6075 ( .A1(net246434), .A2(n4747), .ZN(n4728) );
  NAND2_X2 U6076 ( .A1(n6332), .A2(n6331), .ZN(n6507) );
  NAND2_X4 U6077 ( .A1(n4475), .A2(n4476), .ZN(net245802) );
  NAND2_X2 U6078 ( .A1(n4954), .A2(n4918), .ZN(n4475) );
  INV_X2 U6079 ( .A(n6021), .ZN(n5965) );
  NAND2_X4 U6080 ( .A1(n5925), .A2(n5926), .ZN(n6038) );
  INV_X2 U6081 ( .A(n5958), .ZN(n5957) );
  NAND2_X4 U6082 ( .A1(net245765), .A2(net245764), .ZN(n5065) );
  OAI21_X2 U6083 ( .B1(n3890), .B2(n6611), .A(net243725), .ZN(n6850) );
  INV_X2 U6084 ( .A(n7074), .ZN(n7068) );
  OAI211_X2 U6085 ( .C1(net244278), .C2(n6237), .A(n6236), .B(net244281), .ZN(
        n6238) );
  NOR2_X2 U6086 ( .A1(n7097), .A2(n7096), .ZN(n7101) );
  INV_X2 U6087 ( .A(n6840), .ZN(n6838) );
  NAND2_X2 U6088 ( .A1(n7195), .A2(n4455), .ZN(n7196) );
  XNOR2_X1 U6089 ( .A(n7079), .B(n7078), .ZN(n7010) );
  NAND3_X4 U6090 ( .A1(n4994), .A2(n4992), .A3(n4993), .ZN(n4995) );
  NAND2_X4 U6091 ( .A1(n6069), .A2(n6068), .ZN(n6178) );
  NAND4_X2 U6092 ( .A1(n4839), .A2(n4837), .A3(n4836), .A4(n4835), .ZN(n4886)
         );
  NAND2_X1 U6093 ( .A1(n8025), .A2(n8024), .ZN(n8180) );
  OAI21_X1 U6094 ( .B1(n8025), .B2(n8024), .A(n8023), .ZN(n8181) );
  NOR2_X2 U6095 ( .A1(n4388), .A2(n6771), .ZN(n6775) );
  XNOR2_X2 U6096 ( .A(net245737), .B(net248083), .ZN(n4979) );
  INV_X2 U6097 ( .A(net245737), .ZN(net245739) );
  NAND2_X1 U6098 ( .A1(n6986), .A2(n6985), .ZN(n6801) );
  NAND2_X2 U6099 ( .A1(net247751), .A2(net247752), .ZN(n4505) );
  OAI21_X4 U6100 ( .B1(n4683), .B2(n5294), .A(net245250), .ZN(n4766) );
  NAND2_X2 U6101 ( .A1(net246506), .A2(n4682), .ZN(n4677) );
  NAND2_X4 U6102 ( .A1(net246506), .A2(n4682), .ZN(n4683) );
  NAND2_X2 U6103 ( .A1(n4473), .A2(n4474), .ZN(n4476) );
  INV_X1 U6104 ( .A(n4954), .ZN(n4473) );
  INV_X4 U6105 ( .A(n4918), .ZN(n4474) );
  OAI221_X1 U6106 ( .B1(net246770), .B2(net247083), .C1(net246958), .C2(n6901), 
        .A(n6700), .ZN(n7825) );
  OAI211_X1 U6107 ( .C1(net246770), .C2(n5404), .A(n5403), .B(n5402), .ZN(
        n5432) );
  NOR2_X1 U6108 ( .A1(net246770), .A2(n8298), .ZN(n8299) );
  NAND2_X1 U6109 ( .A1(n5292), .A2(net246770), .ZN(n4599) );
  NAND2_X2 U6110 ( .A1(n7004), .A2(n7003), .ZN(n6843) );
  OAI21_X2 U6111 ( .B1(n7006), .B2(n7005), .A(n7004), .ZN(n7184) );
  NAND2_X4 U6112 ( .A1(n7225), .A2(n7224), .ZN(net242906) );
  NAND2_X2 U6113 ( .A1(n4523), .A2(n4524), .ZN(n6653) );
  OAI21_X4 U6114 ( .B1(net244522), .B2(net244523), .A(n6041), .ZN(n6042) );
  NAND2_X4 U6115 ( .A1(n8538), .A2(n8154), .ZN(n8268) );
  NAND2_X4 U6116 ( .A1(n8094), .A2(n8093), .ZN(n8154) );
  INV_X2 U6117 ( .A(n8085), .ZN(n8087) );
  NAND3_X2 U6118 ( .A1(n7063), .A2(n7073), .A3(n7064), .ZN(n7062) );
  INV_X8 U6119 ( .A(n5129), .ZN(n4509) );
  INV_X8 U6120 ( .A(n4892), .ZN(n5027) );
  NOR3_X4 U6121 ( .A1(n5006), .A2(n5007), .A3(n5005), .ZN(n5026) );
  INV_X4 U6122 ( .A(n8083), .ZN(n8088) );
  NAND2_X4 U6123 ( .A1(n6800), .A2(n6799), .ZN(n6985) );
  OAI21_X2 U6124 ( .B1(n6796), .B2(n6795), .A(n6794), .ZN(n6798) );
  OAI211_X2 U6125 ( .C1(n4006), .C2(net242911), .A(net242908), .B(net242910), 
        .ZN(n7272) );
  NAND3_X1 U6126 ( .A1(net243291), .A2(net243293), .A3(net243294), .ZN(n6936)
         );
  NAND2_X2 U6127 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  OAI21_X4 U6128 ( .B1(n6088), .B2(n6087), .A(n4020), .ZN(n6223) );
  INV_X4 U6129 ( .A(net243311), .ZN(net248038) );
  NAND2_X4 U6130 ( .A1(n6192), .A2(n6191), .ZN(n6358) );
  NAND2_X2 U6131 ( .A1(n5131), .A2(n5130), .ZN(n5133) );
  NAND2_X2 U6132 ( .A1(n6822), .A2(n6826), .ZN(n4482) );
  INV_X8 U6133 ( .A(n7018), .ZN(n7015) );
  NAND2_X2 U6134 ( .A1(net248029), .A2(net248030), .ZN(net248031) );
  XNOR2_X2 U6135 ( .A(n5930), .B(n5929), .ZN(n4478) );
  OAI21_X2 U6136 ( .B1(n6525), .B2(n6660), .A(n6661), .ZN(n6526) );
  NAND2_X2 U6137 ( .A1(n4883), .A2(net245981), .ZN(n4497) );
  NAND2_X2 U6138 ( .A1(n7232), .A2(n7231), .ZN(net242885) );
  OAI21_X1 U6139 ( .B1(n8567), .B2(n8566), .A(n8565), .ZN(n8744) );
  OAI21_X1 U6140 ( .B1(n8571), .B2(n8570), .A(n8569), .ZN(n8742) );
  NOR2_X1 U6141 ( .A1(n8497), .A2(n8498), .ZN(n8501) );
  NAND2_X1 U6142 ( .A1(n8498), .A2(n8497), .ZN(n8499) );
  NAND2_X1 U6143 ( .A1(n7328), .A2(n7327), .ZN(n7133) );
  NAND2_X4 U6144 ( .A1(n5894), .A2(n5893), .ZN(n6075) );
  XNOR2_X2 U6145 ( .A(n6486), .B(n6485), .ZN(n6369) );
  NAND2_X4 U6146 ( .A1(n6810), .A2(n6809), .ZN(n6989) );
  NAND2_X4 U6147 ( .A1(n5076), .A2(n5077), .ZN(n5082) );
  INV_X4 U6148 ( .A(n5078), .ZN(n5076) );
  NAND2_X4 U6149 ( .A1(n4894), .A2(n4893), .ZN(n5004) );
  NAND2_X4 U6150 ( .A1(n6517), .A2(n6516), .ZN(n6655) );
  NAND2_X4 U6151 ( .A1(n6371), .A2(n6370), .ZN(n6494) );
  XNOR2_X2 U6152 ( .A(n5057), .B(n5059), .ZN(n4479) );
  NAND2_X2 U6153 ( .A1(n6222), .A2(n6038), .ZN(n6040) );
  OAI21_X4 U6154 ( .B1(n5136), .B2(n5135), .A(n5134), .ZN(n5915) );
  NAND2_X2 U6155 ( .A1(n4480), .A2(n4481), .ZN(n4483) );
  INV_X1 U6156 ( .A(n6826), .ZN(n4481) );
  NAND2_X4 U6157 ( .A1(a[18]), .A2(b[23]), .ZN(n6826) );
  INV_X8 U6158 ( .A(n6165), .ZN(n6166) );
  NAND2_X4 U6159 ( .A1(n4802), .A2(n4834), .ZN(n4836) );
  NAND2_X4 U6160 ( .A1(n6640), .A2(n6639), .ZN(n6766) );
  NAND2_X4 U6161 ( .A1(n5103), .A2(n5102), .ZN(n5878) );
  INV_X4 U6162 ( .A(n4956), .ZN(n5007) );
  NAND2_X4 U6163 ( .A1(n8042), .A2(n8043), .ZN(n8494) );
  NAND3_X4 U6164 ( .A1(n8041), .A2(n8040), .A3(n8039), .ZN(n8043) );
  NAND2_X4 U6165 ( .A1(n5902), .A2(n5903), .ZN(n6081) );
  NAND2_X4 U6166 ( .A1(n7132), .A2(n7131), .ZN(n7327) );
  INV_X2 U6167 ( .A(n8536), .ZN(n8254) );
  OAI21_X4 U6168 ( .B1(n8171), .B2(n4392), .A(n8169), .ZN(n8507) );
  NAND2_X4 U6169 ( .A1(n4962), .A2(n3956), .ZN(n4994) );
  NAND2_X4 U6170 ( .A1(n8028), .A2(n4432), .ZN(n8029) );
  NAND2_X1 U6171 ( .A1(n7155), .A2(n7154), .ZN(n7156) );
  NOR2_X1 U6172 ( .A1(n7154), .A2(n7155), .ZN(n7158) );
  NAND2_X1 U6173 ( .A1(n6485), .A2(n6486), .ZN(n6488) );
  OAI21_X4 U6174 ( .B1(net244368), .B2(net244369), .A(net244370), .ZN(n6328)
         );
  NOR2_X2 U6175 ( .A1(n8542), .A2(n8541), .ZN(n8545) );
  NAND2_X4 U6176 ( .A1(net241829), .A2(net241824), .ZN(net241756) );
  NOR2_X2 U6177 ( .A1(n6016), .A2(n6015), .ZN(n6019) );
  NAND2_X1 U6178 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  XNOR2_X2 U6179 ( .A(n7389), .B(n4469), .ZN(n7390) );
  NAND2_X2 U6180 ( .A1(n7857), .A2(n7856), .ZN(n4486) );
  NAND2_X4 U6181 ( .A1(n4484), .A2(n4485), .ZN(n4487) );
  NAND2_X4 U6182 ( .A1(n4486), .A2(n4487), .ZN(n7821) );
  INV_X4 U6183 ( .A(n7857), .ZN(n4484) );
  INV_X4 U6184 ( .A(n7856), .ZN(n4485) );
  XNOR2_X2 U6185 ( .A(n7679), .B(net249183), .ZN(n7680) );
  NAND2_X4 U6186 ( .A1(net241751), .A2(n8148), .ZN(n8328) );
  NAND2_X4 U6187 ( .A1(n7682), .A2(n7681), .ZN(net242076) );
  OAI21_X4 U6188 ( .B1(n5016), .B2(n5017), .A(n5015), .ZN(n5023) );
  NAND2_X2 U6189 ( .A1(n6460), .A2(n6461), .ZN(n6621) );
  AOI21_X2 U6190 ( .B1(n3904), .B2(n6097), .A(n4053), .ZN(n5949) );
  NAND2_X4 U6191 ( .A1(n6939), .A2(net243270), .ZN(n6940) );
  NAND2_X2 U6192 ( .A1(n5909), .A2(n5908), .ZN(n4489) );
  NAND2_X4 U6193 ( .A1(n4409), .A2(n4488), .ZN(n4490) );
  NAND2_X4 U6194 ( .A1(n4490), .A2(n4489), .ZN(n5129) );
  NAND2_X4 U6195 ( .A1(a[22]), .A2(b[25]), .ZN(n5908) );
  NAND2_X4 U6196 ( .A1(net246902), .A2(net246768), .ZN(n5452) );
  INV_X8 U6197 ( .A(n4771), .ZN(n4491) );
  INV_X8 U6198 ( .A(n4376), .ZN(n4771) );
  OAI21_X2 U6199 ( .B1(n5901), .B2(n5900), .A(n5899), .ZN(n5904) );
  OAI21_X2 U6200 ( .B1(net246076), .B2(net246075), .A(net248615), .ZN(
        net245910) );
  OAI221_X2 U6201 ( .B1(net244260), .B2(n6240), .C1(net244260), .C2(n6241), 
        .A(n6101), .ZN(n6102) );
  INV_X1 U6202 ( .A(n6822), .ZN(n6824) );
  INV_X2 U6203 ( .A(n5021), .ZN(n5020) );
  OAI21_X2 U6204 ( .B1(net242898), .B2(net242899), .A(net242900), .ZN(
        net242896) );
  NAND2_X4 U6205 ( .A1(n6382), .A2(n6381), .ZN(n6430) );
  OAI21_X4 U6206 ( .B1(net243433), .B2(n6865), .A(n6864), .ZN(n6866) );
  NOR2_X2 U6207 ( .A1(n5014), .A2(n4397), .ZN(n5016) );
  OAI21_X2 U6208 ( .B1(n8166), .B2(n8165), .A(n8164), .ZN(n8517) );
  NOR2_X1 U6209 ( .A1(n7956), .A2(n7957), .ZN(n7960) );
  NAND2_X1 U6210 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  OAI21_X4 U6211 ( .B1(n5049), .B2(net245794), .A(n5048), .ZN(n5053) );
  NAND2_X1 U6212 ( .A1(n6747), .A2(n6746), .ZN(n6749) );
  NAND3_X2 U6213 ( .A1(n6330), .A2(n6329), .A3(n6328), .ZN(n6331) );
  NAND3_X2 U6214 ( .A1(n7887), .A2(n7886), .A3(n7885), .ZN(n7889) );
  NOR2_X2 U6215 ( .A1(n4455), .A2(n7195), .ZN(n7198) );
  INV_X4 U6216 ( .A(n5120), .ZN(n5124) );
  OAI21_X4 U6217 ( .B1(n6162), .B2(n6034), .A(n6160), .ZN(n6035) );
  NAND2_X2 U6218 ( .A1(n7702), .A2(n8071), .ZN(n8072) );
  INV_X2 U6219 ( .A(n8048), .ZN(n8050) );
  NOR2_X2 U6220 ( .A1(n7527), .A2(n7528), .ZN(n7531) );
  NOR2_X2 U6221 ( .A1(n7394), .A2(n7393), .ZN(n7397) );
  NAND2_X4 U6222 ( .A1(n4847), .A2(n4846), .ZN(n4850) );
  XNOR2_X1 U6223 ( .A(n4859), .B(n4815), .ZN(n4769) );
  OAI21_X2 U6224 ( .B1(n4812), .B2(n4815), .A(n4859), .ZN(n4861) );
  NAND2_X4 U6225 ( .A1(a[23]), .A2(net248517), .ZN(n4815) );
  INV_X4 U6226 ( .A(net246070), .ZN(net246076) );
  NAND2_X4 U6227 ( .A1(net249231), .A2(net246754), .ZN(n4767) );
  NAND3_X2 U6228 ( .A1(net246760), .A2(net243754), .A3(net243755), .ZN(n6602)
         );
  NOR2_X2 U6229 ( .A1(n6025), .A2(n6024), .ZN(n6028) );
  NAND2_X4 U6230 ( .A1(n4811), .A2(n4506), .ZN(n4852) );
  NAND2_X4 U6231 ( .A1(n4962), .A2(n4961), .ZN(n4992) );
  XNOR2_X2 U6232 ( .A(net247741), .B(net247843), .ZN(net246576) );
  NAND2_X4 U6233 ( .A1(n5085), .A2(n5084), .ZN(net244674) );
  NAND2_X4 U6234 ( .A1(n4869), .A2(n4870), .ZN(n4912) );
  NAND2_X4 U6235 ( .A1(n6226), .A2(n6225), .ZN(n6230) );
  NAND2_X2 U6236 ( .A1(net246186), .A2(net246105), .ZN(n4492) );
  NAND2_X4 U6237 ( .A1(net247807), .A2(n4492), .ZN(n4880) );
  INV_X4 U6238 ( .A(net246186), .ZN(net247804) );
  NAND2_X2 U6239 ( .A1(net246558), .A2(net246557), .ZN(n4493) );
  NAND2_X4 U6240 ( .A1(net247808), .A2(net247809), .ZN(n4494) );
  NAND2_X4 U6241 ( .A1(n4494), .A2(n4493), .ZN(net245465) );
  INV_X4 U6242 ( .A(net246557), .ZN(net247808) );
  INV_X4 U6243 ( .A(net246558), .ZN(net247809) );
  NAND2_X4 U6244 ( .A1(n4497), .A2(n4498), .ZN(n5439) );
  INV_X1 U6245 ( .A(net245981), .ZN(net247817) );
  NAND2_X1 U6246 ( .A1(net246387), .A2(net248893), .ZN(n4499) );
  NAND2_X4 U6247 ( .A1(n4499), .A2(n4500), .ZN(n4744) );
  INV_X2 U6248 ( .A(net246387), .ZN(net247820) );
  INV_X1 U6249 ( .A(net248717), .ZN(net246558) );
  OAI211_X4 U6250 ( .C1(n4740), .C2(n4744), .A(n4739), .B(n4738), .ZN(
        net246274) );
  NAND2_X2 U6251 ( .A1(n5919), .A2(n5914), .ZN(n4502) );
  NAND2_X4 U6252 ( .A1(n4501), .A2(n5921), .ZN(n4503) );
  NAND2_X2 U6253 ( .A1(n4502), .A2(n4503), .ZN(n5138) );
  INV_X1 U6254 ( .A(n5919), .ZN(n4501) );
  NAND2_X4 U6255 ( .A1(a[23]), .A2(b[24]), .ZN(n5919) );
  NOR2_X1 U6256 ( .A1(n7364), .A2(n7363), .ZN(n7365) );
  NOR2_X1 U6257 ( .A1(n4023), .A2(n6812), .ZN(n6816) );
  NAND2_X1 U6258 ( .A1(n4023), .A2(n6812), .ZN(n6814) );
  NAND2_X4 U6259 ( .A1(n4709), .A2(n4710), .ZN(n4711) );
  XNOR2_X2 U6260 ( .A(n4414), .B(n4920), .ZN(n4923) );
  NAND2_X4 U6261 ( .A1(net246916), .A2(a[30]), .ZN(n4678) );
  NAND2_X4 U6262 ( .A1(b[17]), .A2(a[30]), .ZN(n5954) );
  NAND2_X4 U6263 ( .A1(b[1]), .A2(a[30]), .ZN(n8656) );
  NAND2_X4 U6264 ( .A1(n4803), .A2(n4804), .ZN(n4834) );
  NAND2_X2 U6265 ( .A1(net245808), .A2(n4410), .ZN(n5054) );
  NAND2_X2 U6266 ( .A1(n4415), .A2(n5897), .ZN(n5899) );
  INV_X4 U6267 ( .A(net246384), .ZN(net247762) );
  XNOR2_X2 U6268 ( .A(n4880), .B(n4879), .ZN(n4882) );
  NAND2_X2 U6269 ( .A1(n6384), .A2(n6383), .ZN(net244006) );
  NOR2_X2 U6270 ( .A1(n4740), .A2(n4739), .ZN(n4735) );
  NAND2_X4 U6271 ( .A1(net246327), .A2(n4761), .ZN(n4717) );
  NAND2_X2 U6272 ( .A1(net244665), .A2(net244666), .ZN(n4504) );
  INV_X4 U6273 ( .A(net244666), .ZN(net247752) );
  INV_X8 U6274 ( .A(n5937), .ZN(n6093) );
  INV_X1 U6275 ( .A(net244546), .ZN(net244543) );
  INV_X8 U6276 ( .A(n4893), .ZN(n4958) );
  NAND2_X4 U6277 ( .A1(n4690), .A2(n4689), .ZN(net246385) );
  XNOR2_X2 U6278 ( .A(n5132), .B(n5063), .ZN(net245621) );
  NAND2_X4 U6279 ( .A1(n6241), .A2(n6240), .ZN(net244262) );
  NAND2_X2 U6280 ( .A1(net245786), .A2(net245785), .ZN(n5064) );
  NAND2_X4 U6281 ( .A1(n4867), .A2(n4868), .ZN(net246135) );
  NAND2_X2 U6282 ( .A1(n4699), .A2(n3849), .ZN(n4701) );
  NAND2_X1 U6283 ( .A1(net246760), .A2(b[7]), .ZN(n8758) );
  NAND2_X1 U6284 ( .A1(net246760), .A2(b[8]), .ZN(n8266) );
  AOI22_X1 U6285 ( .A1(n5985), .A2(n4569), .B1(n5449), .B2(net246760), .ZN(
        n5483) );
  XNOR2_X1 U6286 ( .A(net246760), .B(n5309), .ZN(n5310) );
  OAI21_X1 U6287 ( .B1(net248516), .B2(net246762), .A(net245250), .ZN(n5319)
         );
  NOR2_X1 U6288 ( .A1(b[25]), .A2(net246760), .ZN(n5333) );
  OAI221_X1 U6289 ( .B1(net240852), .B2(n8298), .C1(net246958), .C2(net246762), 
        .A(n5162), .ZN(n5787) );
  AOI22_X1 U6290 ( .A1(net247082), .A2(a[17]), .B1(n8834), .B2(net246760), 
        .ZN(n8792) );
  NOR2_X1 U6291 ( .A1(b[25]), .A2(net246762), .ZN(n5505) );
  NAND2_X1 U6292 ( .A1(b[25]), .A2(net246762), .ZN(n5504) );
  NAND2_X1 U6293 ( .A1(net246760), .A2(b[14]), .ZN(n7221) );
  AND2_X2 U6294 ( .A1(n4782), .A2(n4786), .ZN(n4506) );
  INV_X4 U6295 ( .A(n4506), .ZN(n4810) );
  NAND2_X4 U6296 ( .A1(n4775), .A2(n4774), .ZN(n4781) );
  NOR2_X2 U6297 ( .A1(n6973), .A2(n6974), .ZN(n6977) );
  INV_X4 U6298 ( .A(n4747), .ZN(n4748) );
  AND2_X4 U6299 ( .A1(n4781), .A2(n4778), .ZN(n4790) );
  INV_X2 U6300 ( .A(n4778), .ZN(n4782) );
  NAND2_X1 U6301 ( .A1(n4567), .A2(net246754), .ZN(n4778) );
  OAI21_X4 U6302 ( .B1(n6188), .B2(n6187), .A(n6186), .ZN(n6190) );
  NOR2_X4 U6303 ( .A1(net246535), .A2(n4679), .ZN(net246545) );
  NAND2_X4 U6304 ( .A1(net247659), .A2(net247660), .ZN(n4508) );
  NAND2_X4 U6305 ( .A1(n4507), .A2(n4508), .ZN(net245614) );
  INV_X2 U6306 ( .A(net245740), .ZN(net247659) );
  INV_X4 U6307 ( .A(net245741), .ZN(net247660) );
  NAND3_X1 U6308 ( .A1(net243066), .A2(n7078), .A3(net243096), .ZN(n7359) );
  NAND2_X4 U6309 ( .A1(n5127), .A2(n5130), .ZN(n5128) );
  NAND2_X1 U6310 ( .A1(n6982), .A2(n6981), .ZN(n6791) );
  NAND2_X1 U6311 ( .A1(n6358), .A2(n6359), .ZN(n6193) );
  NAND2_X4 U6312 ( .A1(n6492), .A2(n6491), .ZN(n6649) );
  INV_X4 U6313 ( .A(n6490), .ZN(n6492) );
  NAND2_X4 U6314 ( .A1(net246443), .A2(n4708), .ZN(net246345) );
  NAND2_X4 U6315 ( .A1(n4714), .A2(n4777), .ZN(n4756) );
  INV_X4 U6316 ( .A(n6466), .ZN(n6363) );
  NOR2_X4 U6317 ( .A1(n5888), .A2(n5889), .ZN(n5892) );
  NOR2_X2 U6318 ( .A1(n6782), .A2(n6783), .ZN(n6786) );
  NAND2_X1 U6319 ( .A1(net245675), .A2(net245674), .ZN(net245752) );
  NAND4_X2 U6320 ( .A1(net246117), .A2(n4874), .A3(net246118), .A4(net246120), 
        .ZN(net246077) );
  NAND2_X4 U6321 ( .A1(n6743), .A2(n6742), .ZN(n7089) );
  OAI21_X2 U6322 ( .B1(n6741), .B2(n6740), .A(n6739), .ZN(n6742) );
  NAND2_X4 U6323 ( .A1(n6049), .A2(n5913), .ZN(n6039) );
  NAND2_X1 U6324 ( .A1(n6617), .A2(n6616), .ZN(n6474) );
  NOR2_X2 U6325 ( .A1(n6196), .A2(n6197), .ZN(n6200) );
  INV_X2 U6326 ( .A(n4955), .ZN(n4960) );
  NAND2_X4 U6327 ( .A1(n4955), .A2(n5005), .ZN(n4892) );
  INV_X4 U6328 ( .A(net245786), .ZN(net245783) );
  NAND2_X4 U6329 ( .A1(net246578), .A2(net246577), .ZN(net246539) );
  INV_X1 U6330 ( .A(net245988), .ZN(net247630) );
  INV_X2 U6331 ( .A(net247540), .ZN(net245764) );
  NAND3_X2 U6332 ( .A1(n6309), .A2(net244181), .A3(net244180), .ZN(net243775)
         );
  XNOR2_X1 U6333 ( .A(n4904), .B(n4864), .ZN(n4865) );
  NAND2_X4 U6334 ( .A1(n4905), .A2(n4904), .ZN(n4906) );
  OAI21_X2 U6335 ( .B1(n4768), .B2(n3932), .A(n3955), .ZN(n4860) );
  NOR2_X4 U6336 ( .A1(n6890), .A2(n6886), .ZN(n6894) );
  NAND2_X1 U6337 ( .A1(n6153), .A2(n6152), .ZN(n6304) );
  NOR2_X2 U6338 ( .A1(n5897), .A2(n4415), .ZN(n5901) );
  NAND2_X1 U6339 ( .A1(n6849), .A2(n6851), .ZN(n6854) );
  XNOR2_X2 U6340 ( .A(n5133), .B(n5132), .ZN(n5135) );
  NAND2_X1 U6341 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  INV_X2 U6342 ( .A(net244674), .ZN(net245700) );
  NAND2_X4 U6343 ( .A1(n6092), .A2(n3965), .ZN(n6090) );
  NAND2_X4 U6344 ( .A1(n5905), .A2(n5904), .ZN(n6080) );
  OAI21_X4 U6345 ( .B1(n4902), .B2(n4901), .A(n4472), .ZN(n4962) );
  INV_X4 U6346 ( .A(n4568), .ZN(n4567) );
  INV_X2 U6347 ( .A(net244669), .ZN(net245703) );
  NAND2_X1 U6348 ( .A1(n4947), .A2(n4913), .ZN(n4915) );
  INV_X2 U6349 ( .A(n4416), .ZN(n4774) );
  NAND2_X4 U6350 ( .A1(b[31]), .A2(a[29]), .ZN(net246564) );
  NAND2_X2 U6351 ( .A1(n5129), .A2(n5910), .ZN(n4511) );
  NAND2_X4 U6352 ( .A1(n4509), .A2(n4510), .ZN(n4512) );
  NAND2_X4 U6353 ( .A1(n4511), .A2(n4512), .ZN(n5914) );
  INV_X1 U6354 ( .A(n5910), .ZN(n4510) );
  INV_X2 U6355 ( .A(net247549), .ZN(net245711) );
  NAND2_X1 U6356 ( .A1(b[29]), .A2(a[31]), .ZN(net246566) );
  NOR2_X4 U6357 ( .A1(n4401), .A2(n5864), .ZN(n5868) );
  NAND2_X2 U6358 ( .A1(n6456), .A2(n6455), .ZN(n6457) );
  NAND2_X1 U6359 ( .A1(n5915), .A2(n5918), .ZN(n5137) );
  NAND2_X2 U6360 ( .A1(n5918), .A2(n5915), .ZN(n5917) );
  OAI22_X4 U6361 ( .A1(n4960), .A2(n4959), .B1(n5014), .B2(n4397), .ZN(n5033)
         );
  XNOR2_X2 U6362 ( .A(n4479), .B(n5064), .ZN(net247540) );
  OAI21_X1 U6363 ( .B1(n7372), .B2(n4419), .A(n7371), .ZN(n7373) );
  INV_X8 U6364 ( .A(n6885), .ZN(n6890) );
  NAND2_X4 U6365 ( .A1(net243179), .A2(net248987), .ZN(net243106) );
  NAND3_X2 U6366 ( .A1(n8074), .A2(n8073), .A3(n8072), .ZN(n8076) );
  INV_X2 U6367 ( .A(n6866), .ZN(n6869) );
  OAI21_X2 U6368 ( .B1(n6434), .B2(n6433), .A(n6432), .ZN(n6436) );
  NAND2_X4 U6369 ( .A1(n4513), .A2(n4514), .ZN(n4516) );
  NAND2_X4 U6370 ( .A1(n4515), .A2(n4516), .ZN(n7074) );
  INV_X4 U6371 ( .A(n7061), .ZN(n4513) );
  INV_X4 U6372 ( .A(n7060), .ZN(n4514) );
  NAND2_X2 U6373 ( .A1(n7632), .A2(n7633), .ZN(n4519) );
  NAND2_X4 U6374 ( .A1(n4517), .A2(n4518), .ZN(n4520) );
  NAND2_X4 U6375 ( .A1(n4519), .A2(n4520), .ZN(n8082) );
  INV_X4 U6376 ( .A(n7633), .ZN(n4517) );
  INV_X4 U6377 ( .A(n7632), .ZN(n4518) );
  XNOR2_X2 U6378 ( .A(n8082), .B(n7802), .ZN(n7813) );
  NAND2_X1 U6379 ( .A1(n6587), .A2(n6586), .ZN(n6588) );
  NOR2_X2 U6380 ( .A1(n6148), .A2(n6147), .ZN(n6151) );
  NAND2_X1 U6381 ( .A1(net244145), .A2(n6316), .ZN(n6237) );
  NAND2_X4 U6382 ( .A1(net243066), .A2(net243096), .ZN(n7079) );
  NAND2_X4 U6383 ( .A1(n6223), .A2(n6222), .ZN(n6219) );
  NAND2_X4 U6384 ( .A1(n6525), .A2(n6660), .ZN(n6661) );
  NAND2_X4 U6385 ( .A1(n6523), .A2(n6522), .ZN(n6660) );
  INV_X8 U6386 ( .A(net246181), .ZN(net245988) );
  NOR2_X1 U6387 ( .A1(n8518), .A2(n8517), .ZN(n8521) );
  NAND2_X1 U6388 ( .A1(n8518), .A2(n8517), .ZN(n8519) );
  NOR2_X1 U6389 ( .A1(n8508), .A2(n8507), .ZN(n8511) );
  NAND2_X1 U6390 ( .A1(n8508), .A2(n8507), .ZN(n8509) );
  NOR2_X1 U6391 ( .A1(n7987), .A2(n7986), .ZN(n7990) );
  NAND2_X1 U6392 ( .A1(n7987), .A2(n7986), .ZN(n7988) );
  NOR2_X1 U6393 ( .A1(n7976), .A2(n7977), .ZN(n7980) );
  NAND2_X1 U6394 ( .A1(n7977), .A2(n7976), .ZN(n7978) );
  NOR2_X1 U6395 ( .A1(n7936), .A2(n7937), .ZN(n7940) );
  NAND2_X1 U6396 ( .A1(n7937), .A2(n7936), .ZN(n7938) );
  INV_X1 U6397 ( .A(n4899), .ZN(n4521) );
  NAND2_X1 U6398 ( .A1(n6802), .A2(n4522), .ZN(n4523) );
  NAND2_X2 U6399 ( .A1(n4386), .A2(n6803), .ZN(n4524) );
  INV_X4 U6400 ( .A(n6803), .ZN(n4522) );
  OAI21_X2 U6401 ( .B1(n4958), .B2(n4957), .A(n4956), .ZN(n4955) );
  INV_X4 U6402 ( .A(net244659), .ZN(net244655) );
  NAND2_X4 U6403 ( .A1(n4827), .A2(n4828), .ZN(net246100) );
  NAND2_X2 U6404 ( .A1(net246332), .A2(net249177), .ZN(n4698) );
  NAND3_X2 U6405 ( .A1(n4933), .A2(n4934), .A3(n4935), .ZN(n4975) );
  INV_X16 U6406 ( .A(net246918), .ZN(net246916) );
  NAND2_X4 U6407 ( .A1(n4889), .A2(n4413), .ZN(n4893) );
  NAND2_X2 U6408 ( .A1(n5115), .A2(n5113), .ZN(n5024) );
  NAND2_X4 U6409 ( .A1(n6029), .A2(net244535), .ZN(n6161) );
  NAND3_X2 U6410 ( .A1(n6473), .A2(n6472), .A3(n6471), .ZN(n6616) );
  NAND2_X4 U6411 ( .A1(n6600), .A2(n6599), .ZN(net243405) );
  INV_X1 U6412 ( .A(n5370), .ZN(n5371) );
  NAND2_X1 U6413 ( .A1(n7287), .A2(n7286), .ZN(n7595) );
  AND2_X4 U6414 ( .A1(net242602), .A2(n7437), .ZN(n4525) );
  NAND3_X2 U6415 ( .A1(n5023), .A2(n5022), .A3(n5021), .ZN(n5113) );
  NAND2_X4 U6416 ( .A1(n6731), .A2(n6730), .ZN(n6862) );
  INV_X4 U6417 ( .A(n6320), .ZN(n6239) );
  NAND3_X2 U6418 ( .A1(n4949), .A2(n4915), .A3(n4916), .ZN(n4917) );
  NAND2_X4 U6419 ( .A1(n7079), .A2(n7080), .ZN(n7361) );
  NAND2_X4 U6420 ( .A1(n6324), .A2(n6323), .ZN(n6519) );
  NAND2_X1 U6421 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  NAND3_X2 U6422 ( .A1(n4916), .A2(n4915), .A3(n4949), .ZN(n5031) );
  NAND3_X2 U6423 ( .A1(n4491), .A2(n4711), .A3(n4783), .ZN(n4788) );
  NAND3_X4 U6424 ( .A1(n7820), .A2(a[31]), .A3(b[5]), .ZN(n7857) );
  XNOR2_X2 U6425 ( .A(n6363), .B(n6465), .ZN(n6364) );
  NAND2_X2 U6426 ( .A1(n5100), .A2(n5101), .ZN(n5879) );
  XOR2_X1 U6427 ( .A(n6051), .B(n6037), .Z(n4526) );
  XOR2_X2 U6428 ( .A(n6039), .B(n4526), .Z(n5928) );
  NAND2_X4 U6429 ( .A1(b[23]), .A2(a[23]), .ZN(n6037) );
  INV_X4 U6430 ( .A(net248780), .ZN(net243094) );
  AOI21_X1 U6431 ( .B1(n8104), .B2(n7840), .A(n7839), .ZN(n7853) );
  NAND2_X2 U6432 ( .A1(n3954), .A2(n4877), .ZN(n4830) );
  NAND2_X2 U6433 ( .A1(net246188), .A2(n4829), .ZN(n4877) );
  INV_X2 U6434 ( .A(net246342), .ZN(net246434) );
  NOR3_X2 U6435 ( .A1(n7450), .A2(net242581), .A3(net242580), .ZN(n7271) );
  NAND2_X1 U6436 ( .A1(a[30]), .A2(b[4]), .ZN(n8278) );
  NAND3_X1 U6437 ( .A1(a[30]), .A2(n8841), .A3(n1671), .ZN(n5224) );
  OAI21_X1 U6438 ( .B1(net248516), .B2(a[30]), .A(n5236), .ZN(n5748) );
  AOI22_X1 U6439 ( .A1(n4538), .A2(a[31]), .B1(n8318), .B2(a[30]), .ZN(n5248)
         );
  XNOR2_X1 U6440 ( .A(n5231), .B(a[30]), .ZN(n5234) );
  AOI21_X1 U6441 ( .B1(net246962), .B2(a[30]), .A(n6125), .ZN(n5241) );
  AOI22_X1 U6442 ( .A1(net247082), .A2(a[22]), .B1(n8834), .B2(a[30]), .ZN(
        n7420) );
  OAI21_X1 U6443 ( .B1(a[30]), .B2(n5232), .A(n4585), .ZN(n4586) );
  OAI21_X2 U6444 ( .B1(net241746), .B2(n8151), .A(net241493), .ZN(n8152) );
  NAND2_X1 U6445 ( .A1(n8070), .A2(n8071), .ZN(n8074) );
  NAND2_X1 U6446 ( .A1(n7895), .A2(n7894), .ZN(n7899) );
  NAND2_X1 U6447 ( .A1(n7896), .A2(n7894), .ZN(n7898) );
  NOR2_X1 U6448 ( .A1(n7903), .A2(n7902), .ZN(n7906) );
  NAND2_X1 U6449 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  NOR2_X1 U6450 ( .A1(n7967), .A2(n7966), .ZN(n7970) );
  NAND2_X1 U6451 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  NOR2_X1 U6452 ( .A1(n7916), .A2(n7917), .ZN(n7920) );
  NAND2_X1 U6453 ( .A1(n7917), .A2(n7916), .ZN(n7918) );
  NAND2_X1 U6454 ( .A1(n7119), .A2(n7120), .ZN(n7323) );
  NAND2_X4 U6455 ( .A1(net246450), .A2(net248742), .ZN(n4707) );
  NAND2_X1 U6456 ( .A1(n6945), .A2(n6946), .ZN(n6950) );
  NOR2_X2 U6457 ( .A1(n6456), .A2(n6455), .ZN(n6459) );
  XNOR2_X1 U6458 ( .A(n5118), .B(n5864), .ZN(n5885) );
  NOR2_X1 U6459 ( .A1(n5264), .A2(net246776), .ZN(n4596) );
  OAI21_X1 U6460 ( .B1(net248517), .B2(net246776), .A(n5266), .ZN(n5267) );
  OAI221_X1 U6461 ( .B1(net246776), .B2(net247083), .C1(net246958), .C2(n6712), 
        .A(n6565), .ZN(n7658) );
  OAI221_X1 U6462 ( .B1(net245313), .B2(n5378), .C1(net246776), .C2(n5404), 
        .A(n5377), .ZN(n5400) );
  NAND2_X1 U6463 ( .A1(n5264), .A2(net246776), .ZN(n4594) );
  OAI21_X2 U6464 ( .B1(n4954), .B2(n4953), .A(n4952), .ZN(n4972) );
  NAND3_X2 U6465 ( .A1(net246070), .A2(net246072), .A3(net246071), .ZN(n4884)
         );
  AOI21_X4 U6466 ( .B1(n4853), .B2(n4852), .A(n4851), .ZN(n4855) );
  NAND2_X4 U6467 ( .A1(n5039), .A2(n5038), .ZN(n5040) );
  NAND2_X4 U6468 ( .A1(n5089), .A2(n5088), .ZN(n5887) );
  OAI21_X1 U6469 ( .B1(net241491), .B2(net241492), .A(net241493), .ZN(n8338)
         );
  OAI21_X1 U6470 ( .B1(n8540), .B2(n8539), .A(n8538), .ZN(n8541) );
  INV_X2 U6471 ( .A(n4407), .ZN(n8271) );
  INV_X2 U6472 ( .A(n4400), .ZN(n8055) );
  AOI21_X2 U6473 ( .B1(n8053), .B2(n8052), .A(n7705), .ZN(n7778) );
  NAND2_X1 U6474 ( .A1(n7599), .A2(n4465), .ZN(n7588) );
  OAI21_X1 U6475 ( .B1(n4465), .B2(n7599), .A(n7597), .ZN(n7587) );
  INV_X2 U6476 ( .A(n7091), .ZN(n6846) );
  NOR2_X2 U6477 ( .A1(n7090), .A2(n7091), .ZN(n6958) );
  NAND2_X1 U6478 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  NAND2_X4 U6479 ( .A1(n5887), .A2(n5886), .ZN(n5090) );
  OAI211_X4 U6480 ( .C1(n4958), .C2(n4957), .A(n4959), .B(n4956), .ZN(n5002)
         );
  NAND2_X4 U6481 ( .A1(net246016), .A2(net246017), .ZN(n4919) );
  INV_X8 U6482 ( .A(n4919), .ZN(n4927) );
  OAI21_X2 U6483 ( .B1(n5126), .B2(n5125), .A(n4373), .ZN(n5127) );
  NAND2_X4 U6484 ( .A1(n4688), .A2(n4687), .ZN(net246384) );
  NAND2_X4 U6485 ( .A1(n4680), .A2(n5284), .ZN(n4688) );
  NAND2_X4 U6486 ( .A1(n7446), .A2(n7447), .ZN(n8081) );
  OAI21_X2 U6487 ( .B1(n4713), .B2(n4712), .A(n4395), .ZN(n4714) );
  NAND2_X4 U6488 ( .A1(net244541), .A2(net244540), .ZN(n5931) );
  INV_X2 U6489 ( .A(n6883), .ZN(n6595) );
  NAND2_X1 U6490 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  NAND2_X4 U6491 ( .A1(n6728), .A2(n6727), .ZN(n6729) );
  NAND2_X4 U6492 ( .A1(n6942), .A2(n6943), .ZN(net243096) );
  NAND2_X4 U6493 ( .A1(n5266), .A2(n5294), .ZN(net246509) );
  NAND3_X2 U6494 ( .A1(net246289), .A2(net246287), .A3(net246288), .ZN(
        net246238) );
  XNOR2_X2 U6495 ( .A(n4469), .B(n7439), .ZN(n7800) );
  INV_X2 U6496 ( .A(n7876), .ZN(n7682) );
  NAND2_X1 U6497 ( .A1(n8329), .A2(net241503), .ZN(n8331) );
  OAI21_X1 U6498 ( .B1(net241503), .B2(n8329), .A(n3981), .ZN(n8330) );
  NAND2_X1 U6499 ( .A1(n8009), .A2(n8010), .ZN(n8014) );
  NAND3_X1 U6500 ( .A1(n8012), .A2(n8009), .A3(n8011), .ZN(n8015) );
  NAND2_X1 U6501 ( .A1(n4013), .A2(n7184), .ZN(n7186) );
  NOR2_X1 U6502 ( .A1(n7165), .A2(n7164), .ZN(n7168) );
  NAND2_X1 U6503 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  NOR2_X1 U6504 ( .A1(n7135), .A2(n7134), .ZN(n7138) );
  NAND2_X1 U6505 ( .A1(n7135), .A2(n7134), .ZN(n7136) );
  NOR2_X1 U6506 ( .A1(n7125), .A2(n7124), .ZN(n7128) );
  NAND2_X1 U6507 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  NAND2_X1 U6508 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  NOR2_X2 U6509 ( .A1(n6632), .A2(n6633), .ZN(n6636) );
  NOR2_X2 U6510 ( .A1(n6347), .A2(n6348), .ZN(n6351) );
  NOR2_X2 U6511 ( .A1(n6061), .A2(n6062), .ZN(n6065) );
  NOR2_X1 U6512 ( .A1(net241826), .A2(net241749), .ZN(n8101) );
  INV_X2 U6513 ( .A(n8096), .ZN(n8098) );
  NOR2_X2 U6514 ( .A1(n6540), .A2(n6539), .ZN(n6543) );
  NAND2_X1 U6515 ( .A1(net247473), .A2(net241068), .ZN(n8751) );
  INV_X4 U6516 ( .A(n4744), .ZN(n4737) );
  NAND2_X1 U6517 ( .A1(n6388), .A2(n6261), .ZN(n6296) );
  OAI211_X1 U6518 ( .C1(n6388), .C2(net246970), .A(net247048), .B(n6258), .ZN(
        n6259) );
  NAND2_X4 U6519 ( .A1(net245918), .A2(a[24]), .ZN(net245799) );
  NOR2_X2 U6520 ( .A1(n7290), .A2(n7289), .ZN(n7293) );
  NOR2_X4 U6521 ( .A1(n7795), .A2(n8088), .ZN(n7634) );
  INV_X1 U6522 ( .A(n5834), .ZN(n5835) );
  NAND3_X2 U6523 ( .A1(net246497), .A2(net246481), .A3(net246483), .ZN(n4685)
         );
  OAI21_X2 U6524 ( .B1(n7866), .B2(n7862), .A(n7861), .ZN(n7868) );
  NAND2_X4 U6525 ( .A1(n4927), .A2(n4928), .ZN(net245920) );
  INV_X2 U6526 ( .A(net246386), .ZN(net246382) );
  XNOR2_X2 U6527 ( .A(net247847), .B(net244055), .ZN(n6533) );
  NAND3_X1 U6528 ( .A1(n4698), .A2(n4766), .A3(n4716), .ZN(n4699) );
  NAND3_X1 U6529 ( .A1(n5912), .A2(n5911), .A3(n6045), .ZN(n5913) );
  NAND2_X4 U6530 ( .A1(n4715), .A2(n4767), .ZN(n4761) );
  NAND2_X4 U6531 ( .A1(net247778), .A2(net246327), .ZN(n4715) );
  OAI211_X4 U6532 ( .C1(net243759), .C2(net243760), .A(net243757), .B(
        net243761), .ZN(n6601) );
  NAND2_X1 U6533 ( .A1(n7452), .A2(n4468), .ZN(n7453) );
  NOR2_X1 U6534 ( .A1(n7452), .A2(n7573), .ZN(n7454) );
  OAI22_X4 U6535 ( .A1(n5935), .A2(n5934), .B1(n6024), .B2(n6025), .ZN(n5936)
         );
  XNOR2_X2 U6536 ( .A(n6877), .B(n4527), .ZN(n6678) );
  AOI22_X4 U6537 ( .A1(n4807), .A2(n4835), .B1(n4806), .B2(n4805), .ZN(
        net246132) );
  NAND3_X4 U6538 ( .A1(n4837), .A2(n4836), .A3(n4839), .ZN(n4805) );
  XNOR2_X2 U6539 ( .A(n4924), .B(n4945), .ZN(n4928) );
  INV_X1 U6540 ( .A(n4478), .ZN(n6032) );
  INV_X4 U6541 ( .A(net244702), .ZN(net247167) );
  NAND2_X4 U6542 ( .A1(n4790), .A2(n4789), .ZN(n4808) );
  AOI21_X2 U6543 ( .B1(n8763), .B2(net240980), .A(net240981), .ZN(n8765) );
  AOI21_X2 U6544 ( .B1(net244143), .B2(net244144), .A(n6317), .ZN(n6319) );
  NAND2_X4 U6545 ( .A1(net247544), .A2(net244287), .ZN(net244144) );
  NAND2_X1 U6546 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  NOR2_X1 U6547 ( .A1(n7145), .A2(n7144), .ZN(n7148) );
  INV_X1 U6548 ( .A(net246552), .ZN(net245546) );
  OAI21_X4 U6549 ( .B1(n4754), .B2(net246342), .A(n4753), .ZN(n4758) );
  OAI21_X4 U6550 ( .B1(n4748), .B2(net246342), .A(net246353), .ZN(n4749) );
  NAND3_X4 U6551 ( .A1(n4705), .A2(n4704), .A3(n4703), .ZN(net246342) );
  OAI211_X4 U6552 ( .C1(net243866), .C2(net243760), .A(net243761), .B(
        net243757), .ZN(net243781) );
  OAI221_X2 U6553 ( .B1(net246497), .B2(net246483), .C1(net246483), .C2(
        net246481), .A(n4685), .ZN(n4686) );
  XNOR2_X2 U6554 ( .A(net243778), .B(net249128), .ZN(n6598) );
  OAI21_X2 U6555 ( .B1(a[28]), .B2(n5158), .A(n4590), .ZN(n4591) );
  NAND2_X4 U6556 ( .A1(n6087), .A2(n6088), .ZN(n6222) );
  INV_X2 U6557 ( .A(net246908), .ZN(net246904) );
  OAI21_X4 U6558 ( .B1(n6890), .B2(n6891), .A(n6889), .ZN(n6892) );
  OAI21_X2 U6559 ( .B1(n3965), .B2(n6092), .A(n6090), .ZN(n5944) );
  NAND3_X2 U6560 ( .A1(net244260), .A2(n6240), .A3(n6241), .ZN(n6101) );
  NAND2_X4 U6561 ( .A1(n6217), .A2(n6216), .ZN(n6365) );
  OAI21_X2 U6562 ( .B1(n6486), .B2(n6485), .A(n3969), .ZN(n6487) );
  OAI21_X4 U6563 ( .B1(n5075), .B2(n4459), .A(n5073), .ZN(n5078) );
  NAND2_X4 U6564 ( .A1(n7364), .A2(n7363), .ZN(n7083) );
  NAND2_X4 U6565 ( .A1(n6494), .A2(n6495), .ZN(n6496) );
  NAND2_X4 U6566 ( .A1(n6668), .A2(n6667), .ZN(n6748) );
  NAND3_X2 U6567 ( .A1(n6224), .A2(n6223), .A3(n6222), .ZN(n6225) );
  NAND3_X2 U6568 ( .A1(n4728), .A2(net248511), .A3(n4727), .ZN(net246401) );
  NAND2_X1 U6569 ( .A1(n6650), .A2(n6649), .ZN(n6493) );
  INV_X2 U6570 ( .A(n5904), .ZN(n5902) );
  NAND2_X1 U6571 ( .A1(n5122), .A2(n5120), .ZN(n5056) );
  NAND2_X4 U6572 ( .A1(net243271), .A2(n6940), .ZN(n7064) );
  OAI21_X2 U6573 ( .B1(net243433), .B2(n6865), .A(n6864), .ZN(n6878) );
  NOR2_X2 U6574 ( .A1(n5072), .A2(net245722), .ZN(n5075) );
  NAND2_X4 U6575 ( .A1(n4732), .A2(n4743), .ZN(n4738) );
  NAND2_X1 U6576 ( .A1(n4773), .A2(n4772), .ZN(n4783) );
  NAND2_X4 U6577 ( .A1(n4825), .A2(n4824), .ZN(n4875) );
  NAND2_X4 U6578 ( .A1(a[28]), .A2(b[30]), .ZN(n5294) );
  NAND2_X4 U6579 ( .A1(b[29]), .A2(a[30]), .ZN(net245422) );
  NAND2_X4 U6580 ( .A1(n4528), .A2(n4529), .ZN(net245617) );
  NOR2_X4 U6581 ( .A1(n4937), .A2(n4938), .ZN(n4940) );
  NAND2_X4 U6582 ( .A1(net247167), .A2(net247168), .ZN(n4529) );
  NAND2_X4 U6583 ( .A1(net244689), .A2(net244690), .ZN(net245732) );
  NAND2_X4 U6584 ( .A1(n4809), .A2(n4808), .ZN(n4853) );
  NAND2_X2 U6585 ( .A1(net244704), .A2(net244702), .ZN(n4528) );
  INV_X8 U6586 ( .A(n4981), .ZN(n4937) );
  NAND2_X4 U6587 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  NAND2_X4 U6588 ( .A1(n4891), .A2(n4414), .ZN(n4956) );
  NAND2_X4 U6589 ( .A1(n4832), .A2(n4833), .ZN(net246181) );
  NAND2_X4 U6590 ( .A1(n4937), .A2(n4938), .ZN(n4939) );
  NAND2_X4 U6591 ( .A1(n6430), .A2(n6429), .ZN(net244005) );
  NAND2_X4 U6592 ( .A1(n5126), .A2(n5125), .ZN(n5130) );
  NAND2_X4 U6593 ( .A1(n4919), .A2(n4925), .ZN(net245806) );
  NAND2_X4 U6594 ( .A1(n4750), .A2(n4749), .ZN(n4803) );
  NAND2_X4 U6595 ( .A1(net245920), .A2(net245919), .ZN(net245801) );
  NAND2_X1 U6596 ( .A1(n7026), .A2(net242879), .ZN(n7057) );
  OAI211_X1 U6597 ( .C1(net249298), .C2(net246970), .A(net247048), .B(n7023), 
        .ZN(n7024) );
  NAND2_X1 U6598 ( .A1(n6687), .A2(n6551), .ZN(n6583) );
  AOI211_X1 U6599 ( .C1(net246974), .C2(n6692), .A(n6690), .B(n4267), .ZN(
        n6724) );
  OAI211_X1 U6600 ( .C1(n4450), .C2(net240784), .A(net247049), .B(n6548), .ZN(
        n6549) );
  NAND2_X1 U6601 ( .A1(n4447), .A2(n6394), .ZN(n6426) );
  OAI211_X1 U6602 ( .C1(n4447), .C2(net246970), .A(net247048), .B(n6391), .ZN(
        n6392) );
  NAND2_X1 U6603 ( .A1(n6113), .A2(n6255), .ZN(n6144) );
  OAI211_X1 U6604 ( .C1(n6255), .C2(net246970), .A(net247049), .B(n6110), .ZN(
        n6111) );
  NAND2_X1 U6605 ( .A1(n6107), .A2(n5972), .ZN(n6012) );
  OAI211_X1 U6606 ( .C1(n4427), .C2(net246970), .A(net247049), .B(n5969), .ZN(
        n5970) );
  INV_X2 U6607 ( .A(n5294), .ZN(n5295) );
  NAND3_X2 U6608 ( .A1(b[17]), .A2(a[31]), .A3(n5855), .ZN(n5955) );
  OAI21_X2 U6609 ( .B1(n4826), .B2(net246190), .A(n4875), .ZN(n4827) );
  NAND2_X4 U6610 ( .A1(n8267), .A2(n8266), .ZN(net241073) );
  NAND2_X4 U6611 ( .A1(n8265), .A2(n8264), .ZN(net241072) );
  INV_X8 U6612 ( .A(n5061), .ZN(n5126) );
  NAND2_X4 U6613 ( .A1(net244271), .A2(net244272), .ZN(net244076) );
  NAND3_X2 U6614 ( .A1(n8263), .A2(n8262), .A3(n8261), .ZN(n8265) );
  NAND2_X4 U6615 ( .A1(n5924), .A2(n5923), .ZN(n6087) );
  OAI21_X2 U6616 ( .B1(n3933), .B2(n5031), .A(n4952), .ZN(n4918) );
  NAND2_X4 U6617 ( .A1(n4944), .A2(n4943), .ZN(n5066) );
  NAND3_X4 U6618 ( .A1(n4874), .A2(net246117), .A3(net246118), .ZN(net246116)
         );
  NAND2_X4 U6619 ( .A1(net243398), .A2(net243293), .ZN(net243292) );
  NAND3_X2 U6620 ( .A1(n5370), .A2(a[31]), .A3(b[23]), .ZN(n4823) );
  OAI21_X4 U6621 ( .B1(n7876), .B2(n7877), .A(n7875), .ZN(net241599) );
  NOR2_X1 U6622 ( .A1(n4021), .A2(net245318), .ZN(n5376) );
  NAND2_X1 U6623 ( .A1(n8082), .A2(n8081), .ZN(n8085) );
  NAND2_X1 U6624 ( .A1(n8083), .A2(n8081), .ZN(n7802) );
  NAND2_X1 U6625 ( .A1(n4435), .A2(n6835), .ZN(n6841) );
  NOR2_X1 U6626 ( .A1(n6802), .A2(n6803), .ZN(n6806) );
  NAND2_X1 U6627 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  NOR2_X1 U6628 ( .A1(n6793), .A2(n6792), .ZN(n6796) );
  NAND2_X1 U6629 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  NAND2_X1 U6630 ( .A1(n4853), .A2(n4852), .ZN(n4821) );
  NAND2_X1 U6631 ( .A1(n4416), .A2(n4779), .ZN(n4786) );
  OAI21_X1 U6632 ( .B1(n4021), .B2(net246332), .A(n4762), .ZN(n4763) );
  INV_X8 U6633 ( .A(net245317), .ZN(net246327) );
  NAND2_X1 U6634 ( .A1(n7218), .A2(n7217), .ZN(n7220) );
  NAND2_X4 U6635 ( .A1(n6874), .A2(net243423), .ZN(n6881) );
  NAND2_X4 U6636 ( .A1(n4696), .A2(net246475), .ZN(net246445) );
  NAND3_X1 U6637 ( .A1(net249352), .A2(net247545), .A3(a[23]), .ZN(n6236) );
  NAND2_X4 U6638 ( .A1(n8273), .A2(n7859), .ZN(net241012) );
  NAND2_X4 U6639 ( .A1(net246432), .A2(net246433), .ZN(n4751) );
  XNOR2_X2 U6640 ( .A(net248651), .B(n7233), .ZN(n7396) );
  NAND2_X4 U6641 ( .A1(net247847), .A2(n6431), .ZN(net243791) );
  NAND2_X4 U6642 ( .A1(n4681), .A2(net246511), .ZN(n4696) );
  OAI21_X4 U6643 ( .B1(n7445), .B2(n3949), .A(n7444), .ZN(n7448) );
  OAI221_X4 U6644 ( .B1(n6871), .B2(n6870), .C1(n6869), .C2(n6871), .A(n6868), 
        .ZN(n6942) );
  NAND2_X4 U6645 ( .A1(n7448), .A2(n7449), .ZN(n8083) );
  NAND3_X4 U6646 ( .A1(net244072), .A2(net244074), .A3(net244073), .ZN(n6433)
         );
  NAND2_X1 U6647 ( .A1(n7646), .A2(n3911), .ZN(n7677) );
  NAND2_X1 U6648 ( .A1(n7436), .A2(n7406), .ZN(n7434) );
  OAI211_X1 U6649 ( .C1(n7436), .C2(net246970), .A(net247049), .B(n7402), .ZN(
        n7403) );
  NAND2_X1 U6650 ( .A1(n4448), .A2(n7238), .ZN(n7268) );
  OAI211_X1 U6651 ( .C1(n4448), .C2(net246970), .A(net247048), .B(n7235), .ZN(
        n7236) );
  NAND2_X1 U6652 ( .A1(n6935), .A2(n6899), .ZN(n6933) );
  NOR2_X1 U6653 ( .A1(n8768), .A2(n8767), .ZN(n8771) );
  NAND2_X1 U6654 ( .A1(n8768), .A2(n8767), .ZN(n8769) );
  OAI211_X1 U6655 ( .C1(n6935), .C2(net246970), .A(net247049), .B(n6896), .ZN(
        n6897) );
  NAND3_X2 U6656 ( .A1(b[6]), .A2(a[31]), .A3(n7436), .ZN(n7816) );
  NAND2_X4 U6657 ( .A1(n6095), .A2(n6094), .ZN(net244384) );
  NAND2_X4 U6658 ( .A1(net241031), .A2(net241030), .ZN(net240991) );
  NAND2_X4 U6659 ( .A1(n4706), .A2(net245541), .ZN(net246432) );
  XNOR2_X2 U6660 ( .A(n4974), .B(net247658), .ZN(net245888) );
  INV_X2 U6661 ( .A(n6023), .ZN(n6027) );
  NOR2_X1 U6662 ( .A1(net240783), .A2(net246970), .ZN(n8860) );
  NAND2_X1 U6663 ( .A1(n4426), .A2(n8286), .ZN(n8325) );
  AOI21_X1 U6664 ( .B1(n8280), .B2(n8129), .A(n8128), .ZN(n8142) );
  NAND2_X1 U6665 ( .A1(n7374), .A2(n7375), .ZN(n7378) );
  NAND2_X1 U6666 ( .A1(n7376), .A2(n7375), .ZN(n7377) );
  NAND3_X1 U6667 ( .A1(n7360), .A2(n7361), .A3(n7363), .ZN(n7367) );
  NAND2_X4 U6668 ( .A1(net243747), .A2(net248442), .ZN(n6728) );
  NAND3_X1 U6669 ( .A1(net249194), .A2(net243734), .A3(net243733), .ZN(n6610)
         );
  NAND2_X1 U6670 ( .A1(n6434), .A2(n6433), .ZN(n6435) );
  INV_X2 U6671 ( .A(n6433), .ZN(n6377) );
  NAND3_X1 U6672 ( .A1(net244143), .A2(net244144), .A3(a[23]), .ZN(n6318) );
  NAND2_X1 U6673 ( .A1(net244545), .A2(n4478), .ZN(n6029) );
  NAND3_X1 U6674 ( .A1(net244540), .A2(net244541), .A3(n4478), .ZN(n6030) );
  NAND3_X2 U6675 ( .A1(net246345), .A2(net246346), .A3(n4751), .ZN(n4747) );
  NAND3_X2 U6676 ( .A1(n4751), .A2(net246346), .A3(net246345), .ZN(n4752) );
  NAND2_X4 U6677 ( .A1(ALUCtrl[2]), .A2(net246918), .ZN(n8312) );
  INV_X16 U6678 ( .A(n4531), .ZN(n8842) );
  INV_X8 U6679 ( .A(n8298), .ZN(n8834) );
  INV_X32 U6680 ( .A(n4532), .ZN(n4533) );
  NAND2_X4 U6681 ( .A1(b[29]), .A2(net246908), .ZN(n8832) );
  NAND2_X4 U6682 ( .A1(ALUCtrl[2]), .A2(net249231), .ZN(n8806) );
  INV_X16 U6683 ( .A(n4535), .ZN(n8125) );
  NAND2_X4 U6684 ( .A1(net245052), .A2(net246920), .ZN(n8848) );
  INV_X16 U6685 ( .A(n4537), .ZN(n8318) );
  NAND2_X4 U6686 ( .A1(net246916), .A2(net245052), .ZN(n8804) );
  INV_X16 U6687 ( .A(n4539), .ZN(n8841) );
  INV_X32 U6688 ( .A(net247059), .ZN(net247060) );
  NAND2_X4 U6689 ( .A1(net246589), .A2(net246932), .ZN(net240917) );
  INV_X16 U6690 ( .A(net247060), .ZN(net240913) );
  INV_X32 U6691 ( .A(n4540), .ZN(n4541) );
  NAND2_X4 U6692 ( .A1(n5150), .A2(net246932), .ZN(n8850) );
  INV_X16 U6693 ( .A(n4541), .ZN(n8784) );
  INV_X32 U6694 ( .A(net241814), .ZN(net247043) );
  INV_X32 U6695 ( .A(net247043), .ZN(net247044) );
  INV_X32 U6696 ( .A(n4544), .ZN(n4542) );
  INV_X32 U6697 ( .A(n4544), .ZN(n4543) );
  INV_X32 U6698 ( .A(n4548), .ZN(n4546) );
  INV_X32 U6699 ( .A(n4548), .ZN(n4547) );
  INV_X32 U6700 ( .A(n4545), .ZN(n4548) );
  INV_X32 U6701 ( .A(n3931), .ZN(n4550) );
  INV_X32 U6702 ( .A(net247048), .ZN(net247002) );
  INV_X32 U6703 ( .A(n4556), .ZN(n4554) );
  INV_X32 U6704 ( .A(n4560), .ZN(n4557) );
  INV_X32 U6705 ( .A(n4560), .ZN(n4558) );
  INV_X32 U6706 ( .A(n4533), .ZN(n4561) );
  INV_X32 U6707 ( .A(net246966), .ZN(net246960) );
  INV_X32 U6708 ( .A(net246966), .ZN(net246962) );
  INV_X32 U6709 ( .A(net246960), .ZN(net246956) );
  INV_X32 U6710 ( .A(net246960), .ZN(net246958) );
  INV_X32 U6711 ( .A(n4563), .ZN(n4564) );
  INV_X32 U6712 ( .A(n4563), .ZN(n4565) );
  INV_X32 U6713 ( .A(n4564), .ZN(n4566) );
  INV_X32 U6714 ( .A(net246930), .ZN(net246924) );
  INV_X32 U6715 ( .A(net246930), .ZN(net246926) );
  INV_X32 U6716 ( .A(ALUCtrl[0]), .ZN(net246930) );
  INV_X32 U6717 ( .A(b[30]), .ZN(net246908) );
  INV_X32 U6718 ( .A(b[29]), .ZN(n4569) );
  INV_X32 U6719 ( .A(net246888), .ZN(net246880) );
  INV_X32 U6720 ( .A(a[30]), .ZN(net246804) );
  INV_X32 U6721 ( .A(net246756), .ZN(net246754) );
  INV_X32 U6722 ( .A(a[21]), .ZN(n4572) );
  INV_X32 U6723 ( .A(a[19]), .ZN(n4575) );
  INV_X32 U6724 ( .A(a[18]), .ZN(n4576) );
  INV_X32 U6725 ( .A(a[17]), .ZN(n4577) );
  INV_X32 U6726 ( .A(n4579), .ZN(n4578) );
  INV_X32 U6727 ( .A(a[16]), .ZN(n4579) );
  INV_X32 U6728 ( .A(a[15]), .ZN(n4580) );
  INV_X32 U6729 ( .A(a[14]), .ZN(n4581) );
  NAND2_X2 U6730 ( .A1(ALUCtrl[3]), .A2(a[0]), .ZN(n8786) );
  INV_X4 U6731 ( .A(n8786), .ZN(n8845) );
  NAND2_X2 U6732 ( .A1(net246958), .A2(n8845), .ZN(n7044) );
  INV_X4 U6733 ( .A(n7044), .ZN(n24) );
  NAND2_X2 U6734 ( .A1(ALUCtrl[3]), .A2(net245052), .ZN(n4669) );
  INV_X4 U6735 ( .A(n4669), .ZN(n4582) );
  NAND2_X2 U6736 ( .A1(ALUCtrl[1]), .A2(n4582), .ZN(n8856) );
  INV_X4 U6737 ( .A(n8856), .ZN(n8781) );
  XNOR2_X2 U6738 ( .A(net246924), .B(b[16]), .ZN(n5975) );
  XNOR2_X2 U6739 ( .A(a[16]), .B(n5975), .ZN(n4627) );
  XNOR2_X2 U6740 ( .A(net246924), .B(b[29]), .ZN(n5204) );
  XNOR2_X2 U6741 ( .A(ALUCtrl[0]), .B(b[31]), .ZN(n5805) );
  NAND2_X2 U6742 ( .A1(net246924), .A2(a[31]), .ZN(n4584) );
  NOR2_X4 U6743 ( .A1(net246924), .A2(a[31]), .ZN(n4583) );
  AOI21_X4 U6744 ( .B1(n5805), .B2(n4584), .A(n4583), .ZN(n5232) );
  NAND2_X2 U6745 ( .A1(n5232), .A2(a[30]), .ZN(n4587) );
  XNOR2_X2 U6746 ( .A(net246926), .B(net246902), .ZN(n5231) );
  INV_X4 U6747 ( .A(n5231), .ZN(n4585) );
  NAND2_X2 U6748 ( .A1(n4587), .A2(n4586), .ZN(n5205) );
  NAND2_X2 U6749 ( .A1(net246786), .A2(n5205), .ZN(n4589) );
  NOR2_X4 U6750 ( .A1(net246790), .A2(n5205), .ZN(n4588) );
  AOI21_X4 U6751 ( .B1(n5204), .B2(n4589), .A(n4588), .ZN(n5158) );
  NAND2_X2 U6752 ( .A1(n5158), .A2(a[28]), .ZN(n4592) );
  XNOR2_X2 U6753 ( .A(net246924), .B(net246878), .ZN(n5156) );
  INV_X4 U6754 ( .A(n5156), .ZN(n4590) );
  NAND2_X2 U6755 ( .A1(n4592), .A2(n4591), .ZN(n4593) );
  INV_X4 U6756 ( .A(n4593), .ZN(n5264) );
  XNOR2_X2 U6757 ( .A(net246924), .B(b[27]), .ZN(n5265) );
  INV_X4 U6758 ( .A(n5265), .ZN(n4595) );
  OAI21_X4 U6759 ( .B1(n4596), .B2(n4595), .A(n4594), .ZN(n5292) );
  XNOR2_X2 U6760 ( .A(net246924), .B(b[26]), .ZN(n5293) );
  INV_X4 U6761 ( .A(n5293), .ZN(n4598) );
  INV_X4 U6762 ( .A(n5292), .ZN(n4597) );
  AOI22_X2 U6763 ( .A1(n4599), .A2(n4598), .B1(n4597), .B2(net246766), .ZN(
        n5311) );
  NOR2_X4 U6764 ( .A1(n5311), .A2(net246762), .ZN(n4602) );
  XNOR2_X2 U6765 ( .A(net246926), .B(b[25]), .ZN(n5309) );
  INV_X4 U6766 ( .A(n5309), .ZN(n4601) );
  NAND2_X2 U6767 ( .A1(n5311), .A2(net246764), .ZN(n4600) );
  OAI21_X4 U6768 ( .B1(n4602), .B2(n4601), .A(n4600), .ZN(n5348) );
  NAND2_X2 U6769 ( .A1(n5348), .A2(net246756), .ZN(n4605) );
  XNOR2_X2 U6770 ( .A(net246926), .B(b[24]), .ZN(n5349) );
  INV_X4 U6771 ( .A(n5349), .ZN(n4604) );
  INV_X4 U6772 ( .A(n5348), .ZN(n4603) );
  AOI22_X2 U6773 ( .A1(n4605), .A2(n4604), .B1(n4603), .B2(a[24]), .ZN(n5365)
         );
  XNOR2_X2 U6774 ( .A(net246926), .B(b[23]), .ZN(n5363) );
  INV_X4 U6775 ( .A(n5363), .ZN(n4607) );
  NAND2_X2 U6776 ( .A1(n5365), .A2(net246750), .ZN(n4606) );
  OAI21_X4 U6777 ( .B1(n4608), .B2(n4607), .A(n4606), .ZN(n5393) );
  NAND2_X2 U6778 ( .A1(n5393), .A2(n4571), .ZN(n4611) );
  XNOR2_X2 U6779 ( .A(net246926), .B(b[22]), .ZN(n5392) );
  INV_X4 U6780 ( .A(n5392), .ZN(n4610) );
  INV_X4 U6781 ( .A(n5393), .ZN(n4609) );
  AOI22_X2 U6782 ( .A1(n4611), .A2(n4610), .B1(n4609), .B2(a[22]), .ZN(n5422)
         );
  XNOR2_X2 U6783 ( .A(net246926), .B(net246836), .ZN(n5423) );
  INV_X4 U6784 ( .A(n5423), .ZN(n4613) );
  NAND2_X2 U6785 ( .A1(n5422), .A2(n4573), .ZN(n4612) );
  OAI21_X4 U6786 ( .B1(n4614), .B2(n4613), .A(n4612), .ZN(n5447) );
  NAND2_X2 U6787 ( .A1(n5447), .A2(n4574), .ZN(n4617) );
  XNOR2_X2 U6788 ( .A(net246926), .B(b[20]), .ZN(n5448) );
  INV_X4 U6789 ( .A(n5448), .ZN(n4616) );
  INV_X4 U6790 ( .A(n5447), .ZN(n4615) );
  AOI22_X2 U6791 ( .A1(n4617), .A2(n4616), .B1(n4615), .B2(a[20]), .ZN(n5472)
         );
  XNOR2_X2 U6792 ( .A(net246926), .B(b[19]), .ZN(n5473) );
  INV_X4 U6793 ( .A(n5473), .ZN(n4619) );
  NAND2_X2 U6794 ( .A1(n5472), .A2(n4575), .ZN(n4618) );
  OAI21_X4 U6795 ( .B1(n4620), .B2(n4619), .A(n4618), .ZN(n5816) );
  NAND2_X2 U6796 ( .A1(n5816), .A2(n4576), .ZN(n4623) );
  XNOR2_X2 U6797 ( .A(net246926), .B(b[18]), .ZN(n5815) );
  INV_X4 U6798 ( .A(n5815), .ZN(n4622) );
  INV_X4 U6799 ( .A(n5816), .ZN(n4621) );
  AOI22_X2 U6800 ( .A1(n4623), .A2(n4622), .B1(n4621), .B2(a[18]), .ZN(n5845)
         );
  XNOR2_X2 U6801 ( .A(net246926), .B(b[17]), .ZN(n5843) );
  INV_X4 U6802 ( .A(n5843), .ZN(n4625) );
  NAND2_X2 U6803 ( .A1(n5845), .A2(n4577), .ZN(n4624) );
  OAI21_X4 U6804 ( .B1(n4626), .B2(n4625), .A(n4624), .ZN(n5976) );
  XNOR2_X2 U6805 ( .A(n4627), .B(n5976), .ZN(n4674) );
  NAND2_X2 U6806 ( .A1(b[27]), .A2(net246878), .ZN(n8298) );
  NAND2_X2 U6807 ( .A1(n8834), .A2(n8845), .ZN(n5314) );
  NAND2_X2 U6808 ( .A1(net246878), .A2(net246876), .ZN(n4628) );
  INV_X4 U6809 ( .A(n4628), .ZN(n5995) );
  NAND2_X2 U6810 ( .A1(n4543), .A2(a[8]), .ZN(n8836) );
  INV_X4 U6811 ( .A(n8836), .ZN(n4630) );
  INV_X4 U6812 ( .A(a[0]), .ZN(net240839) );
  NOR2_X4 U6813 ( .A1(n4630), .A2(n4629), .ZN(n4631) );
  OAI211_X2 U6814 ( .C1(net246958), .C2(n4579), .A(n5314), .B(n4631), .ZN(
        n5474) );
  NAND2_X2 U6815 ( .A1(n5474), .A2(n4565), .ZN(n4640) );
  NAND2_X2 U6816 ( .A1(net246902), .A2(n4569), .ZN(n8115) );
  NOR2_X4 U6817 ( .A1(n8786), .A2(net246874), .ZN(n4645) );
  AOI21_X4 U6818 ( .B1(n4542), .B2(a[6]), .A(n4645), .ZN(n4633) );
  NAND2_X2 U6819 ( .A1(net246962), .A2(a[14]), .ZN(n4632) );
  NAND2_X2 U6820 ( .A1(n4633), .A2(n4632), .ZN(n5994) );
  NAND2_X2 U6821 ( .A1(n4555), .A2(n5994), .ZN(n4639) );
  AOI21_X4 U6822 ( .B1(n4542), .B2(a[2]), .A(n4645), .ZN(n4635) );
  NAND2_X2 U6823 ( .A1(net246962), .A2(a[10]), .ZN(n4634) );
  NAND2_X2 U6824 ( .A1(n4635), .A2(n4634), .ZN(n6560) );
  NAND2_X2 U6825 ( .A1(n4562), .A2(n6560), .ZN(n4638) );
  INV_X4 U6826 ( .A(n8832), .ZN(n8796) );
  NAND2_X2 U6827 ( .A1(net246962), .A2(a[12]), .ZN(n6410) );
  INV_X4 U6828 ( .A(n4645), .ZN(n5997) );
  NAND2_X2 U6829 ( .A1(n4542), .A2(a[4]), .ZN(n4636) );
  NAND3_X2 U6830 ( .A1(n6410), .A2(n5997), .A3(n4636), .ZN(n6273) );
  NAND2_X2 U6831 ( .A1(n4558), .A2(n6273), .ZN(n4637) );
  NAND4_X2 U6832 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n5849)
         );
  AOI21_X4 U6833 ( .B1(n4542), .B2(a[7]), .A(n4645), .ZN(n4642) );
  NAND2_X2 U6834 ( .A1(net246962), .A2(a[15]), .ZN(n4641) );
  NAND2_X2 U6835 ( .A1(n4642), .A2(n4641), .ZN(n5824) );
  NAND2_X2 U6836 ( .A1(n5824), .A2(n4565), .ZN(n4651) );
  NAND2_X2 U6837 ( .A1(net246962), .A2(a[13]), .ZN(n6282) );
  NAND2_X2 U6838 ( .A1(n4542), .A2(a[5]), .ZN(n4643) );
  NAND3_X2 U6839 ( .A1(n6282), .A2(n5997), .A3(n4643), .ZN(n6129) );
  NAND2_X2 U6840 ( .A1(n4555), .A2(n6129), .ZN(n4650) );
  NAND2_X2 U6841 ( .A1(net246962), .A2(a[9]), .ZN(n6918) );
  NAND2_X2 U6842 ( .A1(n4542), .A2(a[1]), .ZN(n4644) );
  NAND3_X2 U6843 ( .A1(n6918), .A2(n5997), .A3(n4644), .ZN(n6697) );
  NAND2_X2 U6844 ( .A1(n4561), .A2(n6697), .ZN(n4649) );
  AOI21_X4 U6845 ( .B1(n4542), .B2(a[3]), .A(n4645), .ZN(n4647) );
  NAND2_X2 U6846 ( .A1(net246962), .A2(a[11]), .ZN(n4646) );
  NAND2_X2 U6847 ( .A1(n4647), .A2(n4646), .ZN(n6404) );
  NAND2_X2 U6848 ( .A1(n4558), .A2(n6404), .ZN(n4648) );
  NAND4_X2 U6849 ( .A1(n4651), .A2(n4650), .A3(n4649), .A4(n4648), .ZN(n5982)
         );
  AOI22_X2 U6850 ( .A1(n8842), .A2(n5849), .B1(n8125), .B2(n5982), .ZN(n4672)
         );
  NAND2_X2 U6851 ( .A1(n4542), .A2(a[30]), .ZN(n4652) );
  OAI21_X4 U6852 ( .B1(net246956), .B2(n4571), .A(n4652), .ZN(n5818) );
  NAND2_X2 U6853 ( .A1(net246962), .A2(a[20]), .ZN(n4654) );
  NAND2_X2 U6854 ( .A1(n4542), .A2(a[28]), .ZN(n4653) );
  NAND2_X2 U6855 ( .A1(n4654), .A2(n4653), .ZN(n5450) );
  INV_X4 U6856 ( .A(n5450), .ZN(n6122) );
  NAND2_X2 U6857 ( .A1(n4542), .A2(net246766), .ZN(n4656) );
  OAI21_X4 U6858 ( .B1(net246956), .B2(n4576), .A(n4656), .ZN(n6408) );
  NAND2_X2 U6859 ( .A1(net246962), .A2(n4578), .ZN(n4658) );
  NAND2_X2 U6860 ( .A1(n4542), .A2(net246754), .ZN(n4657) );
  NAND2_X2 U6861 ( .A1(n4658), .A2(n4657), .ZN(n6699) );
  AOI22_X2 U6862 ( .A1(n4555), .A2(n6408), .B1(n6699), .B2(n4564), .ZN(n4659)
         );
  NAND2_X2 U6863 ( .A1(n4660), .A2(n4659), .ZN(n5981) );
  NAND2_X2 U6864 ( .A1(net246962), .A2(a[21]), .ZN(n4662) );
  NAND2_X2 U6865 ( .A1(n4542), .A2(net246790), .ZN(n4661) );
  NAND2_X2 U6866 ( .A1(n4662), .A2(n4661), .ZN(n5985) );
  NAND2_X2 U6867 ( .A1(n4542), .A2(a[31]), .ZN(n4663) );
  OAI21_X4 U6868 ( .B1(net246956), .B2(net246750), .A(n4663), .ZN(n5480) );
  AOI22_X2 U6869 ( .A1(n5985), .A2(n4559), .B1(n4561), .B2(n5480), .ZN(n4668)
         );
  NAND2_X2 U6870 ( .A1(net246962), .A2(a[17]), .ZN(n4665) );
  NAND2_X2 U6871 ( .A1(n4542), .A2(net246760), .ZN(n4664) );
  NAND2_X2 U6872 ( .A1(n4665), .A2(n4664), .ZN(n6563) );
  NAND2_X2 U6873 ( .A1(n4542), .A2(net246772), .ZN(n4666) );
  OAI21_X4 U6874 ( .B1(net246956), .B2(n4575), .A(n4666), .ZN(n6280) );
  AOI22_X2 U6875 ( .A1(n6563), .A2(n4564), .B1(n4554), .B2(n6280), .ZN(n4667)
         );
  NAND2_X2 U6876 ( .A1(n4668), .A2(n4667), .ZN(n5848) );
  AOI22_X2 U6877 ( .A1(n8318), .A2(n5981), .B1(n8841), .B2(n5848), .ZN(n4671)
         );
  AOI21_X2 U6878 ( .B1(n4552), .B2(n4674), .A(n4673), .ZN(n5155) );
  INV_X4 U6879 ( .A(b[16]), .ZN(net244627) );
  INV_X4 U6880 ( .A(net244867), .ZN(net246589) );
  NOR2_X4 U6881 ( .A1(n4551), .A2(n4675), .ZN(n5149) );
  NAND2_X2 U6882 ( .A1(b[20]), .A2(net246786), .ZN(n4943) );
  INV_X4 U6883 ( .A(n4943), .ZN(n4941) );
  INV_X4 U6884 ( .A(n4983), .ZN(n4938) );
  NOR2_X4 U6885 ( .A1(net247632), .A2(net246868), .ZN(n4680) );
  XOR2_X2 U6886 ( .A(net246534), .B(net245313), .Z(net246569) );
  NAND2_X2 U6887 ( .A1(a[30]), .A2(a[31]), .ZN(n4676) );
  INV_X4 U6888 ( .A(n4677), .ZN(n4679) );
  NAND2_X2 U6889 ( .A1(b[30]), .A2(a[29]), .ZN(n5266) );
  INV_X4 U6890 ( .A(net245313), .ZN(net245393) );
  NOR3_X4 U6891 ( .A1(net246542), .A2(net245393), .A3(net246536), .ZN(
        net246514) );
  NAND2_X2 U6892 ( .A1(b[26]), .A2(a[30]), .ZN(n4687) );
  OAI211_X2 U6893 ( .C1(net246514), .C2(net246513), .A(net245349), .B(
        net246515), .ZN(n4681) );
  NAND2_X2 U6894 ( .A1(n4567), .A2(net246772), .ZN(n4695) );
  XNOR2_X2 U6895 ( .A(n5452), .B(net246463), .ZN(n4691) );
  XNOR2_X2 U6896 ( .A(n4691), .B(n4695), .ZN(n4684) );
  NAND2_X2 U6897 ( .A1(net246878), .A2(net246778), .ZN(net245541) );
  NAND2_X2 U6898 ( .A1(b[27]), .A2(net246786), .ZN(net246483) );
  XNOR2_X2 U6899 ( .A(n4686), .B(net249142), .ZN(net246386) );
  INV_X4 U6900 ( .A(n4687), .ZN(n4690) );
  INV_X4 U6901 ( .A(n4688), .ZN(n4689) );
  NAND2_X2 U6902 ( .A1(net246878), .A2(net246772), .ZN(net246346) );
  XNOR2_X2 U6903 ( .A(n4692), .B(n4691), .ZN(n4697) );
  INV_X4 U6904 ( .A(n4697), .ZN(n4693) );
  INV_X4 U6905 ( .A(n4695), .ZN(n4710) );
  NAND3_X2 U6906 ( .A1(n4697), .A2(n4696), .A3(net246466), .ZN(n4709) );
  XNOR2_X2 U6907 ( .A(n4701), .B(n4700), .ZN(n4772) );
  NAND2_X2 U6908 ( .A1(n4567), .A2(net246768), .ZN(n4784) );
  INV_X4 U6909 ( .A(n4784), .ZN(n4773) );
  NAND3_X2 U6910 ( .A1(n4491), .A2(n4711), .A3(n4106), .ZN(n4705) );
  NAND2_X2 U6911 ( .A1(n4713), .A2(n4702), .ZN(n4704) );
  NAND2_X2 U6912 ( .A1(n4771), .A2(n4702), .ZN(n4703) );
  NAND3_X4 U6913 ( .A1(net246447), .A2(net246448), .A3(n4707), .ZN(net246433)
         );
  INV_X4 U6914 ( .A(net245541), .ZN(net246443) );
  XNOR2_X2 U6915 ( .A(net246445), .B(net248354), .ZN(n4708) );
  INV_X4 U6916 ( .A(net246432), .ZN(net246431) );
  OAI21_X4 U6917 ( .B1(n4713), .B2(n4771), .A(n4773), .ZN(n4777) );
  NOR3_X4 U6918 ( .A1(n4721), .A2(n4720), .A3(n4719), .ZN(n4722) );
  NAND2_X2 U6919 ( .A1(a[23]), .A2(net246916), .ZN(n4764) );
  XNOR2_X2 U6920 ( .A(n4722), .B(n4764), .ZN(n4724) );
  NAND2_X2 U6921 ( .A1(net246904), .A2(net246754), .ZN(n4765) );
  INV_X4 U6922 ( .A(n4765), .ZN(n4723) );
  XNOR2_X2 U6923 ( .A(n4724), .B(n4723), .ZN(n4780) );
  NAND2_X2 U6924 ( .A1(net246760), .A2(n4567), .ZN(n4779) );
  XNOR2_X2 U6925 ( .A(n4780), .B(n4779), .ZN(n4755) );
  INV_X4 U6926 ( .A(n4755), .ZN(n4725) );
  NAND2_X2 U6927 ( .A1(net246878), .A2(net246768), .ZN(n4753) );
  INV_X4 U6928 ( .A(n4753), .ZN(n4750) );
  XNOR2_X2 U6929 ( .A(n4725), .B(n4750), .ZN(n4726) );
  INV_X4 U6930 ( .A(n4729), .ZN(n4727) );
  INV_X4 U6931 ( .A(n4728), .ZN(n4730) );
  NAND2_X2 U6932 ( .A1(net246397), .A2(net246395), .ZN(net246289) );
  XNOR2_X2 U6933 ( .A(net246392), .B(net246393), .ZN(net246273) );
  AOI21_X2 U6934 ( .B1(net246385), .B2(net246386), .A(net247762), .ZN(
        net246389) );
  NAND2_X2 U6935 ( .A1(b[25]), .A2(a[30]), .ZN(n4742) );
  INV_X4 U6936 ( .A(n4742), .ZN(n4732) );
  NAND2_X2 U6937 ( .A1(net246384), .A2(net246385), .ZN(n4731) );
  XNOR2_X2 U6938 ( .A(net246382), .B(n4731), .ZN(n5331) );
  INV_X4 U6939 ( .A(n4733), .ZN(n4743) );
  INV_X4 U6940 ( .A(n4738), .ZN(n4736) );
  NAND2_X2 U6941 ( .A1(n4733), .A2(n4742), .ZN(n4734) );
  INV_X4 U6942 ( .A(n4734), .ZN(n4740) );
  NAND2_X2 U6943 ( .A1(b[25]), .A2(net246786), .ZN(n4739) );
  OAI21_X4 U6944 ( .B1(n4737), .B2(n4736), .A(n4735), .ZN(net246272) );
  XNOR2_X2 U6945 ( .A(net246273), .B(n4741), .ZN(n4800) );
  XNOR2_X2 U6946 ( .A(n4743), .B(n4742), .ZN(n4745) );
  XNOR2_X2 U6947 ( .A(n4745), .B(n4744), .ZN(n5340) );
  XNOR2_X2 U6948 ( .A(n4800), .B(n4798), .ZN(n4746) );
  NAND2_X2 U6949 ( .A1(b[24]), .A2(a[30]), .ZN(n4797) );
  XNOR2_X2 U6950 ( .A(n4746), .B(n4797), .ZN(n5370) );
  NAND2_X2 U6951 ( .A1(net246760), .A2(net246882), .ZN(n4840) );
  INV_X4 U6952 ( .A(net246349), .ZN(net246348) );
  NOR2_X4 U6953 ( .A1(net246346), .A2(net246348), .ZN(n4759) );
  INV_X4 U6954 ( .A(n4752), .ZN(n4754) );
  XNOR2_X2 U6955 ( .A(n4756), .B(n4412), .ZN(n4757) );
  OAI21_X4 U6956 ( .B1(n4758), .B2(n4759), .A(n4757), .ZN(n4804) );
  XNOR2_X2 U6957 ( .A(n4760), .B(n4840), .ZN(n4794) );
  INV_X4 U6958 ( .A(n4860), .ZN(n4816) );
  NOR2_X4 U6959 ( .A1(n4812), .A2(n4816), .ZN(n4770) );
  NAND2_X2 U6960 ( .A1(a[22]), .A2(net249231), .ZN(n4859) );
  XNOR2_X2 U6961 ( .A(n4770), .B(n4769), .ZN(n4809) );
  INV_X4 U6962 ( .A(n4779), .ZN(n4775) );
  NAND4_X2 U6963 ( .A1(n4777), .A2(n4776), .A3(n4781), .A4(n4783), .ZN(n4811)
         );
  NAND3_X2 U6964 ( .A1(n4788), .A2(n4787), .A3(n4786), .ZN(n4789) );
  XNOR2_X2 U6965 ( .A(n4809), .B(n4792), .ZN(n4838) );
  NAND2_X2 U6966 ( .A1(b[27]), .A2(net246768), .ZN(net246239) );
  INV_X4 U6967 ( .A(n4797), .ZN(n4796) );
  INV_X4 U6968 ( .A(n4798), .ZN(n4795) );
  NAND2_X2 U6969 ( .A1(n4796), .A2(n4795), .ZN(net246205) );
  NAND2_X2 U6970 ( .A1(n4798), .A2(n4797), .ZN(n4799) );
  NAND2_X2 U6971 ( .A1(b[24]), .A2(net246786), .ZN(net246204) );
  NAND3_X4 U6972 ( .A1(b[22]), .A2(a[31]), .A3(n5411), .ZN(n4879) );
  NAND2_X2 U6973 ( .A1(b[22]), .A2(a[30]), .ZN(n4881) );
  NAND2_X2 U6974 ( .A1(b[25]), .A2(net246772), .ZN(net246120) );
  XNOR2_X2 U6975 ( .A(net246254), .B(n3930), .ZN(n4801) );
  NAND2_X2 U6976 ( .A1(b[26]), .A2(net246768), .ZN(net245429) );
  INV_X4 U6977 ( .A(net246239), .ZN(net246130) );
  NAND2_X2 U6978 ( .A1(net246130), .A2(net246129), .ZN(n4868) );
  NAND2_X2 U6979 ( .A1(net246760), .A2(b[27]), .ZN(net246127) );
  INV_X4 U6980 ( .A(n4840), .ZN(n4802) );
  NAND2_X2 U6981 ( .A1(n4802), .A2(n4838), .ZN(n4837) );
  NAND2_X2 U6982 ( .A1(net246878), .A2(net246754), .ZN(n4835) );
  INV_X4 U6983 ( .A(n4835), .ZN(n4806) );
  INV_X4 U6984 ( .A(n4861), .ZN(n4814) );
  NAND2_X2 U6985 ( .A1(a[22]), .A2(net248517), .ZN(n4813) );
  NAND2_X2 U6986 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  NAND3_X2 U6987 ( .A1(n4861), .A2(n4817), .A3(a[22]), .ZN(n4863) );
  NAND2_X2 U6988 ( .A1(n4818), .A2(n4863), .ZN(n4843) );
  NAND2_X2 U6989 ( .A1(a[23]), .A2(n4567), .ZN(n4846) );
  NAND2_X2 U6990 ( .A1(a[21]), .A2(net249231), .ZN(n4842) );
  XNOR2_X2 U6991 ( .A(n4846), .B(n4842), .ZN(n4819) );
  XNOR2_X2 U6992 ( .A(n4843), .B(n4819), .ZN(n4820) );
  XNOR2_X2 U6993 ( .A(n4821), .B(n4820), .ZN(net246172) );
  XNOR2_X2 U6994 ( .A(net246003), .B(net246198), .ZN(net246105) );
  INV_X4 U6995 ( .A(n4876), .ZN(n4828) );
  NAND2_X2 U6996 ( .A1(n4823), .A2(n4822), .ZN(n4829) );
  INV_X4 U6997 ( .A(n4829), .ZN(n4826) );
  INV_X4 U6998 ( .A(n4822), .ZN(n4825) );
  INV_X4 U6999 ( .A(n4880), .ZN(n4831) );
  AOI21_X4 U7000 ( .B1(n4879), .B2(n4881), .A(n4831), .ZN(net245989) );
  INV_X4 U7001 ( .A(n4881), .ZN(n4833) );
  NAND2_X2 U7002 ( .A1(b[25]), .A2(net246768), .ZN(net246074) );
  NAND3_X2 U7003 ( .A1(net245429), .A2(net246177), .A3(net246176), .ZN(
        net246179) );
  INV_X4 U7004 ( .A(net246172), .ZN(net246133) );
  NAND2_X2 U7005 ( .A1(net246133), .A2(n4835), .ZN(n4887) );
  NAND3_X2 U7006 ( .A1(n4887), .A2(n4886), .A3(n4885), .ZN(n4920) );
  NAND2_X2 U7007 ( .A1(a[22]), .A2(n4567), .ZN(n4896) );
  INV_X4 U7008 ( .A(n4896), .ZN(n4854) );
  INV_X4 U7009 ( .A(n4846), .ZN(n4845) );
  XNOR2_X2 U7010 ( .A(n4843), .B(n4842), .ZN(n4847) );
  INV_X4 U7011 ( .A(n4847), .ZN(n4844) );
  NAND2_X2 U7012 ( .A1(n4845), .A2(n4844), .ZN(n4897) );
  INV_X4 U7013 ( .A(n4897), .ZN(n4856) );
  NOR2_X4 U7014 ( .A1(n4854), .A2(n4856), .ZN(n4858) );
  INV_X4 U7015 ( .A(n4853), .ZN(n4848) );
  OAI21_X4 U7016 ( .B1(n4849), .B2(n4848), .A(n4850), .ZN(n4895) );
  INV_X4 U7017 ( .A(n4850), .ZN(n4851) );
  OAI21_X4 U7018 ( .B1(n4855), .B2(n4856), .A(n4854), .ZN(n4900) );
  INV_X4 U7019 ( .A(n4900), .ZN(n4857) );
  NAND2_X2 U7020 ( .A1(a[21]), .A2(net246902), .ZN(n4903) );
  NAND3_X2 U7021 ( .A1(n4861), .A2(n4860), .A3(a[21]), .ZN(n4862) );
  NAND3_X2 U7022 ( .A1(n3953), .A2(n4863), .A3(n4862), .ZN(n4904) );
  NAND2_X2 U7023 ( .A1(a[20]), .A2(net246916), .ZN(n4967) );
  XNOR2_X2 U7024 ( .A(n4903), .B(n4967), .ZN(n4864) );
  INV_X4 U7025 ( .A(n4865), .ZN(n4902) );
  XNOR2_X2 U7026 ( .A(n4888), .B(n4902), .ZN(n4921) );
  NAND2_X2 U7027 ( .A1(a[23]), .A2(net246882), .ZN(n4957) );
  XNOR2_X2 U7028 ( .A(n4921), .B(n4957), .ZN(n4866) );
  XNOR2_X2 U7029 ( .A(n4866), .B(n4920), .ZN(n4913) );
  INV_X4 U7030 ( .A(n4913), .ZN(n4872) );
  NAND2_X2 U7031 ( .A1(net246760), .A2(b[26]), .ZN(net245921) );
  NAND2_X2 U7032 ( .A1(b[27]), .A2(net246754), .ZN(n4950) );
  XOR2_X2 U7033 ( .A(net245921), .B(n4950), .Z(n4871) );
  XNOR2_X2 U7034 ( .A(net246132), .B(net246133), .ZN(n4870) );
  NAND3_X2 U7035 ( .A1(n4868), .A2(net246127), .A3(n4867), .ZN(n4869) );
  FA_X1 U7036 ( .A(n4872), .B(n4871), .CI(n4945), .S(n4873) );
  XNOR2_X2 U7037 ( .A(n4873), .B(n4919), .ZN(net246073) );
  XNOR2_X2 U7038 ( .A(net246106), .B(net246107), .ZN(net246086) );
  XNOR2_X2 U7039 ( .A(net246096), .B(net245985), .ZN(n4929) );
  XNOR2_X2 U7040 ( .A(n4882), .B(n4881), .ZN(net245268) );
  INV_X4 U7041 ( .A(net245268), .ZN(net246091) );
  NAND3_X4 U7042 ( .A1(n5439), .A2(a[31]), .A3(b[20]), .ZN(n4981) );
  NAND2_X2 U7043 ( .A1(b[23]), .A2(net246772), .ZN(net246082) );
  INV_X4 U7044 ( .A(net246074), .ZN(net246068) );
  NAND2_X2 U7045 ( .A1(net246068), .A2(n4884), .ZN(net245911) );
  NAND2_X2 U7046 ( .A1(b[25]), .A2(net246760), .ZN(net245369) );
  NAND2_X2 U7047 ( .A1(a[22]), .A2(net246880), .ZN(n4959) );
  INV_X4 U7048 ( .A(n4959), .ZN(n5005) );
  NAND3_X2 U7049 ( .A1(n4887), .A2(n4886), .A3(n4885), .ZN(n4889) );
  INV_X4 U7050 ( .A(n4889), .ZN(n4891) );
  INV_X4 U7051 ( .A(n4957), .ZN(n4894) );
  NAND2_X2 U7052 ( .A1(n4897), .A2(n4896), .ZN(n4898) );
  INV_X4 U7053 ( .A(n4903), .ZN(n4905) );
  NOR2_X4 U7054 ( .A1(n4905), .A2(n4904), .ZN(n4907) );
  OAI21_X4 U7055 ( .B1(n4907), .B2(n4967), .A(n4906), .ZN(n4965) );
  NAND2_X2 U7056 ( .A1(a[20]), .A2(net248516), .ZN(n4964) );
  NAND2_X2 U7057 ( .A1(a[19]), .A2(net246916), .ZN(n4963) );
  XNOR2_X2 U7058 ( .A(n4964), .B(n4963), .ZN(n4908) );
  XNOR2_X2 U7059 ( .A(n4965), .B(n4908), .ZN(n4961) );
  XNOR2_X2 U7060 ( .A(n4909), .B(n4961), .ZN(n4910) );
  XNOR2_X2 U7061 ( .A(n4910), .B(n3956), .ZN(n5028) );
  INV_X4 U7062 ( .A(n5028), .ZN(n5003) );
  XNOR2_X2 U7063 ( .A(n4911), .B(n5003), .ZN(n4954) );
  INV_X4 U7064 ( .A(n4912), .ZN(n4914) );
  INV_X4 U7065 ( .A(net246034), .ZN(net246031) );
  INV_X4 U7066 ( .A(n4950), .ZN(n4947) );
  OAI21_X4 U7067 ( .B1(n4914), .B2(net246031), .A(n4947), .ZN(n4916) );
  XNOR2_X2 U7068 ( .A(n4866), .B(n4920), .ZN(n4946) );
  OAI21_X4 U7069 ( .B1(n4914), .B2(net246031), .A(n4946), .ZN(n4949) );
  NAND2_X2 U7070 ( .A1(n3933), .A2(n4917), .ZN(n4952) );
  XNOR2_X2 U7071 ( .A(n4950), .B(n4957), .ZN(n4922) );
  XNOR2_X2 U7072 ( .A(n4923), .B(n4922), .ZN(n4924) );
  NAND2_X2 U7073 ( .A1(b[26]), .A2(net246754), .ZN(net245805) );
  INV_X4 U7074 ( .A(net246017), .ZN(net246013) );
  OAI21_X4 U7075 ( .B1(net246013), .B2(net246014), .A(n4925), .ZN(n4926) );
  XNOR2_X2 U7076 ( .A(net245991), .B(net245992), .ZN(net245963) );
  XNOR2_X2 U7077 ( .A(net245984), .B(net249300), .ZN(n4977) );
  NAND2_X2 U7078 ( .A1(n3966), .A2(net245981), .ZN(n4934) );
  INV_X4 U7079 ( .A(n4934), .ZN(n4932) );
  NAND2_X2 U7080 ( .A1(net246836), .A2(net246786), .ZN(n4935) );
  INV_X4 U7081 ( .A(n4935), .ZN(n4930) );
  OAI21_X4 U7082 ( .B1(n4932), .B2(n4931), .A(n4930), .ZN(n4976) );
  XNOR2_X2 U7083 ( .A(n4936), .B(n4977), .ZN(n4982) );
  OAI21_X4 U7084 ( .B1(n4940), .B2(n4982), .A(n4939), .ZN(n4942) );
  INV_X4 U7085 ( .A(n4942), .ZN(n4944) );
  AOI21_X2 U7086 ( .B1(n4947), .B2(n4946), .A(n3933), .ZN(n4948) );
  NAND2_X2 U7087 ( .A1(n3956), .A2(n4961), .ZN(n4993) );
  INV_X4 U7088 ( .A(n4995), .ZN(n4998) );
  NAND2_X2 U7089 ( .A1(a[20]), .A2(n4567), .ZN(n4997) );
  INV_X4 U7090 ( .A(n4997), .ZN(n4996) );
  NAND2_X2 U7091 ( .A1(a[19]), .A2(net246902), .ZN(n4988) );
  NAND2_X2 U7092 ( .A1(n4964), .A2(n4963), .ZN(n4966) );
  NAND2_X2 U7093 ( .A1(n4966), .A2(n4965), .ZN(n4987) );
  OAI21_X4 U7094 ( .B1(n4967), .B2(n4988), .A(n4987), .ZN(n4985) );
  NAND2_X2 U7095 ( .A1(a[18]), .A2(net249231), .ZN(n5107) );
  XNOR2_X2 U7096 ( .A(n4988), .B(n5107), .ZN(n4968) );
  XNOR2_X2 U7097 ( .A(n4985), .B(n4968), .ZN(n5008) );
  NAND2_X2 U7098 ( .A1(a[21]), .A2(net246880), .ZN(n5001) );
  XNOR2_X2 U7099 ( .A(n5008), .B(n5001), .ZN(n4969) );
  NAND2_X2 U7100 ( .A1(a[22]), .A2(b[27]), .ZN(n5034) );
  XNOR2_X2 U7101 ( .A(n5032), .B(n5034), .ZN(n4970) );
  XNOR2_X2 U7102 ( .A(n5033), .B(n4970), .ZN(n4971) );
  XNOR2_X2 U7103 ( .A(n4972), .B(n4971), .ZN(n5045) );
  INV_X4 U7104 ( .A(n5045), .ZN(n5046) );
  NAND2_X2 U7105 ( .A1(a[23]), .A2(b[26]), .ZN(n5047) );
  XNOR2_X2 U7106 ( .A(n5046), .B(n5047), .ZN(n4973) );
  INV_X4 U7107 ( .A(net245921), .ZN(net245919) );
  NAND3_X4 U7108 ( .A1(net245805), .A2(net245806), .A3(net245801), .ZN(
        net245810) );
  XNOR2_X2 U7109 ( .A(net245808), .B(n4973), .ZN(n5057) );
  NAND2_X2 U7110 ( .A1(b[25]), .A2(a[24]), .ZN(n5059) );
  INV_X4 U7111 ( .A(net245369), .ZN(net245907) );
  XNOR2_X2 U7112 ( .A(n4479), .B(n5064), .ZN(net245906) );
  NAND2_X2 U7113 ( .A1(net246760), .A2(b[24]), .ZN(net245762) );
  INV_X4 U7114 ( .A(net245888), .ZN(net244689) );
  INV_X4 U7115 ( .A(n4975), .ZN(n4978) );
  OAI21_X4 U7116 ( .B1(n4977), .B2(n4978), .A(n4976), .ZN(net245737) );
  XNOR2_X2 U7117 ( .A(n4979), .B(net244689), .ZN(n5067) );
  XNOR2_X2 U7118 ( .A(n4980), .B(n5069), .ZN(n5074) );
  NAND2_X2 U7119 ( .A1(b[19]), .A2(a[30]), .ZN(n5071) );
  XNOR2_X2 U7120 ( .A(n5074), .B(n5071), .ZN(n4984) );
  XNOR2_X2 U7121 ( .A(n4984), .B(net245722), .ZN(n5834) );
  NAND3_X4 U7122 ( .A1(n5834), .A2(a[31]), .A3(b[18]), .ZN(n5141) );
  NAND2_X2 U7123 ( .A1(b[18]), .A2(a[30]), .ZN(n5140) );
  XOR2_X2 U7124 ( .A(n5141), .B(n5140), .Z(n5081) );
  INV_X4 U7125 ( .A(n4985), .ZN(n4986) );
  NOR2_X4 U7126 ( .A1(n4988), .A2(n4986), .ZN(n4990) );
  NOR2_X4 U7127 ( .A1(n4990), .A2(n4989), .ZN(n5104) );
  NAND2_X2 U7128 ( .A1(a[17]), .A2(net246916), .ZN(n5105) );
  XOR2_X2 U7129 ( .A(n5104), .B(n5105), .Z(n4991) );
  NAND2_X2 U7130 ( .A1(a[18]), .A2(net248516), .ZN(n5106) );
  XNOR2_X2 U7131 ( .A(n4991), .B(n5106), .ZN(n5095) );
  INV_X4 U7132 ( .A(n5008), .ZN(n5092) );
  NAND2_X2 U7133 ( .A1(n4996), .A2(n4995), .ZN(n5091) );
  NAND2_X2 U7134 ( .A1(n5092), .A2(n5091), .ZN(n5096) );
  XNOR2_X2 U7135 ( .A(n4430), .B(n4999), .ZN(n5000) );
  NAND2_X2 U7136 ( .A1(a[19]), .A2(n4567), .ZN(n5098) );
  XNOR2_X2 U7137 ( .A(n5000), .B(n5098), .ZN(n5114) );
  INV_X4 U7138 ( .A(n5001), .ZN(n5012) );
  NAND2_X2 U7139 ( .A1(n5003), .A2(n5002), .ZN(n5010) );
  OAI21_X4 U7140 ( .B1(n5007), .B2(n5006), .A(n5005), .ZN(n5013) );
  NAND3_X2 U7141 ( .A1(n5010), .A2(n5013), .A3(n4396), .ZN(n5011) );
  INV_X4 U7142 ( .A(n5013), .ZN(n5017) );
  INV_X4 U7143 ( .A(n5023), .ZN(n5019) );
  NAND2_X2 U7144 ( .A1(a[20]), .A2(net246880), .ZN(n5022) );
  INV_X4 U7145 ( .A(n5022), .ZN(n5018) );
  OAI21_X4 U7146 ( .B1(n5020), .B2(n5019), .A(n5018), .ZN(n5115) );
  XNOR2_X2 U7147 ( .A(n5114), .B(n5024), .ZN(n5089) );
  NAND2_X2 U7148 ( .A1(a[21]), .A2(b[27]), .ZN(n5025) );
  INV_X4 U7149 ( .A(n5025), .ZN(n5041) );
  XNOR2_X2 U7150 ( .A(n4911), .B(n4397), .ZN(n5030) );
  XNOR2_X2 U7151 ( .A(n5033), .B(n5032), .ZN(n5035) );
  AOI21_X4 U7152 ( .B1(n5037), .B2(n5036), .A(n5035), .ZN(n5042) );
  INV_X4 U7153 ( .A(n5034), .ZN(n5039) );
  NAND3_X2 U7154 ( .A1(n5037), .A2(n5036), .A3(n5035), .ZN(n5038) );
  INV_X4 U7155 ( .A(n5040), .ZN(n5043) );
  OAI21_X4 U7156 ( .B1(n5043), .B2(n5042), .A(n5041), .ZN(n5886) );
  INV_X4 U7157 ( .A(n5054), .ZN(n5052) );
  INV_X4 U7158 ( .A(net245806), .ZN(net245803) );
  INV_X4 U7159 ( .A(net245805), .ZN(net245804) );
  NAND2_X2 U7160 ( .A1(n5046), .A2(net245799), .ZN(n5049) );
  INV_X4 U7161 ( .A(n5047), .ZN(n5048) );
  INV_X4 U7162 ( .A(n5053), .ZN(n5051) );
  NAND2_X2 U7163 ( .A1(a[22]), .A2(b[26]), .ZN(n5055) );
  INV_X4 U7164 ( .A(n5055), .ZN(n5050) );
  OAI21_X4 U7165 ( .B1(n5052), .B2(n5051), .A(n5050), .ZN(n5122) );
  NAND3_X2 U7166 ( .A1(n5055), .A2(n5054), .A3(n5053), .ZN(n5120) );
  INV_X4 U7167 ( .A(net245785), .ZN(net245782) );
  OAI21_X4 U7168 ( .B1(n5060), .B2(n5059), .A(n5058), .ZN(n5061) );
  NAND2_X2 U7169 ( .A1(a[23]), .A2(b[25]), .ZN(n5125) );
  INV_X4 U7170 ( .A(n5125), .ZN(n5062) );
  NAND2_X2 U7171 ( .A1(n5130), .A2(n5131), .ZN(n5063) );
  INV_X4 U7172 ( .A(net245768), .ZN(net245761) );
  OAI21_X4 U7173 ( .B1(net245761), .B2(net245762), .A(n5065), .ZN(n5134) );
  NAND2_X2 U7174 ( .A1(b[24]), .A2(a[24]), .ZN(n5345) );
  XNOR2_X2 U7175 ( .A(n5134), .B(n5345), .ZN(net245760) );
  NAND2_X2 U7176 ( .A1(net246836), .A2(net246772), .ZN(net244688) );
  NAND2_X2 U7177 ( .A1(net245732), .A2(net245731), .ZN(net245615) );
  INV_X4 U7178 ( .A(n5066), .ZN(n5070) );
  INV_X4 U7179 ( .A(n5067), .ZN(n5069) );
  XNOR2_X2 U7180 ( .A(n5085), .B(n5086), .ZN(net245724) );
  INV_X4 U7181 ( .A(n5071), .ZN(n5072) );
  NAND2_X2 U7182 ( .A1(n5072), .A2(net245722), .ZN(n5073) );
  NAND2_X2 U7183 ( .A1(b[19]), .A2(net246786), .ZN(n5077) );
  XNOR2_X2 U7184 ( .A(net245711), .B(n5080), .ZN(n5145) );
  XNOR2_X2 U7185 ( .A(n5081), .B(n5145), .ZN(n5855) );
  INV_X4 U7186 ( .A(n5955), .ZN(n5951) );
  XNOR2_X2 U7187 ( .A(n5951), .B(n5954), .ZN(n5148) );
  NAND2_X2 U7188 ( .A1(b[19]), .A2(a[28]), .ZN(n5938) );
  XNOR2_X2 U7189 ( .A(n5938), .B(n5083), .ZN(n5139) );
  INV_X4 U7190 ( .A(n5086), .ZN(n5084) );
  NAND2_X2 U7191 ( .A1(b[20]), .A2(net246772), .ZN(net244567) );
  INV_X4 U7192 ( .A(net244567), .ZN(net245698) );
  NAND2_X2 U7193 ( .A1(b[23]), .A2(a[24]), .ZN(net244704) );
  NAND2_X2 U7194 ( .A1(a[20]), .A2(b[27]), .ZN(n5891) );
  XNOR2_X2 U7195 ( .A(n5090), .B(n5891), .ZN(n5119) );
  NAND2_X2 U7196 ( .A1(a[18]), .A2(n4567), .ZN(n5102) );
  INV_X4 U7197 ( .A(n5102), .ZN(n5100) );
  NAND2_X2 U7198 ( .A1(n5092), .A2(n5091), .ZN(n5093) );
  NAND3_X2 U7199 ( .A1(n5096), .A2(n5095), .A3(n5094), .ZN(n5097) );
  INV_X4 U7200 ( .A(n5101), .ZN(n5103) );
  NAND2_X2 U7201 ( .A1(n5879), .A2(n5878), .ZN(n5112) );
  NAND2_X2 U7202 ( .A1(a[17]), .A2(net248517), .ZN(n5872) );
  NOR2_X4 U7203 ( .A1(n5109), .A2(n5108), .ZN(n5873) );
  INV_X4 U7204 ( .A(n5873), .ZN(n5111) );
  NAND2_X2 U7205 ( .A1(n4578), .A2(net249231), .ZN(n5871) );
  XNOR2_X2 U7206 ( .A(n5872), .B(n5871), .ZN(n5110) );
  XNOR2_X2 U7207 ( .A(n5111), .B(n5110), .ZN(n5877) );
  XNOR2_X2 U7208 ( .A(n5112), .B(n5877), .ZN(n5865) );
  NAND2_X2 U7209 ( .A1(a[19]), .A2(net246880), .ZN(n5867) );
  XNOR2_X2 U7210 ( .A(n5865), .B(n5867), .ZN(n5118) );
  INV_X4 U7211 ( .A(n5113), .ZN(n5117) );
  INV_X4 U7212 ( .A(n5114), .ZN(n5116) );
  OAI21_X4 U7213 ( .B1(n5117), .B2(n5116), .A(n5115), .ZN(n5864) );
  XNOR2_X2 U7214 ( .A(n5119), .B(n4420), .ZN(n5898) );
  OAI21_X4 U7215 ( .B1(n5124), .B2(n5123), .A(n5122), .ZN(n5897) );
  NAND2_X2 U7216 ( .A1(a[21]), .A2(b[26]), .ZN(n5900) );
  INV_X4 U7217 ( .A(n5345), .ZN(n5136) );
  NAND2_X2 U7218 ( .A1(n5136), .A2(net245621), .ZN(n5918) );
  XNOR2_X2 U7219 ( .A(n5138), .B(n5137), .ZN(net244701) );
  INV_X4 U7220 ( .A(n5140), .ZN(n5143) );
  INV_X4 U7221 ( .A(n5141), .ZN(n5142) );
  NAND2_X2 U7222 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  OAI21_X4 U7223 ( .B1(n5146), .B2(n5145), .A(n5144), .ZN(n5945) );
  INV_X4 U7224 ( .A(n5947), .ZN(n5946) );
  OAI22_X2 U7225 ( .A1(n5948), .A2(n5947), .B1(n5946), .B2(n5945), .ZN(n5147)
         );
  XNOR2_X2 U7226 ( .A(n3904), .B(n5147), .ZN(n5958) );
  XNOR2_X2 U7227 ( .A(n5148), .B(n5958), .ZN(n5966) );
  MUX2_X2 U7228 ( .A(n3999), .B(n5149), .S(n4421), .Z(n5154) );
  NAND2_X2 U7229 ( .A1(a[16]), .A2(b[16]), .ZN(n8729) );
  NAND2_X2 U7230 ( .A1(n3991), .A2(n8729), .ZN(n5571) );
  INV_X4 U7231 ( .A(n5571), .ZN(n5152) );
  INV_X4 U7232 ( .A(ALUCtrl[3]), .ZN(net244933) );
  NAND3_X4 U7233 ( .A1(ALUCtrl[2]), .A2(net244841), .A3(net244933), .ZN(n5778)
         );
  INV_X4 U7234 ( .A(n5778), .ZN(n5150) );
  NAND3_X4 U7235 ( .A1(net244841), .A2(net246932), .A3(net245052), .ZN(
        net241814) );
  AOI221_X2 U7236 ( .B1(n5152), .B2(n8784), .C1(n4267), .C2(n3991), .A(n5151), 
        .ZN(n5153) );
  NAND3_X2 U7237 ( .A1(n5155), .A2(n5154), .A3(n5153), .ZN(out[16]) );
  XNOR2_X2 U7238 ( .A(n5156), .B(net246782), .ZN(n5157) );
  XNOR2_X2 U7239 ( .A(n5158), .B(n5157), .ZN(n5159) );
  NAND2_X2 U7240 ( .A1(n8781), .A2(n5159), .ZN(n5203) );
  INV_X4 U7241 ( .A(a[1]), .ZN(net240852) );
  NAND2_X2 U7242 ( .A1(n4543), .A2(a[17]), .ZN(n6919) );
  INV_X4 U7243 ( .A(n6919), .ZN(n5161) );
  INV_X4 U7244 ( .A(a[9]), .ZN(n7029) );
  NOR2_X4 U7245 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  NAND2_X2 U7246 ( .A1(n4555), .A2(n5787), .ZN(n5174) );
  INV_X4 U7247 ( .A(a[5]), .ZN(n7842) );
  NAND2_X2 U7248 ( .A1(n4543), .A2(a[13]), .ZN(n7660) );
  INV_X4 U7249 ( .A(n7660), .ZN(n5163) );
  INV_X4 U7250 ( .A(n5314), .ZN(n5351) );
  NOR2_X4 U7251 ( .A1(n5163), .A2(n5351), .ZN(n5164) );
  OAI221_X2 U7252 ( .B1(n7842), .B2(net247083), .C1(net246958), .C2(n4572), 
        .A(n5164), .ZN(n5395) );
  NAND2_X2 U7253 ( .A1(n4561), .A2(n5395), .ZN(n5173) );
  NAND2_X2 U7254 ( .A1(n4543), .A2(a[15]), .ZN(n7249) );
  NAND2_X2 U7255 ( .A1(net246962), .A2(a[23]), .ZN(n5166) );
  NAND2_X2 U7256 ( .A1(net247082), .A2(a[7]), .ZN(n5165) );
  NAND4_X2 U7257 ( .A1(n5314), .A2(n7249), .A3(n5166), .A4(n5165), .ZN(n5353)
         );
  NAND2_X2 U7258 ( .A1(n4543), .A2(a[19]), .ZN(n6565) );
  INV_X4 U7259 ( .A(n6565), .ZN(n5168) );
  INV_X4 U7260 ( .A(a[11]), .ZN(n6712) );
  NOR2_X4 U7261 ( .A1(n6712), .A2(net247083), .ZN(n5167) );
  NOR2_X4 U7262 ( .A1(n5168), .A2(n5167), .ZN(n5171) );
  INV_X4 U7263 ( .A(a[3]), .ZN(n8289) );
  AOI21_X4 U7264 ( .B1(net246962), .B2(net246772), .A(n5169), .ZN(n5170) );
  NAND2_X2 U7265 ( .A1(n5171), .A2(n5170), .ZN(n5788) );
  AOI22_X2 U7266 ( .A1(n4557), .A2(n5353), .B1(n5788), .B2(n4564), .ZN(n5172)
         );
  NAND3_X2 U7267 ( .A1(n5174), .A2(n5173), .A3(n5172), .ZN(n5277) );
  INV_X4 U7268 ( .A(n5277), .ZN(n5176) );
  NAND2_X2 U7269 ( .A1(net246962), .A2(n4569), .ZN(net245318) );
  NAND2_X2 U7270 ( .A1(net248517), .A2(a[31]), .ZN(net245388) );
  OAI22_X2 U7271 ( .A1(net245318), .A2(net245388), .B1(n620), .B2(net246792), 
        .ZN(n5212) );
  NAND2_X2 U7272 ( .A1(n8841), .A2(n5212), .ZN(n5175) );
  OAI21_X4 U7273 ( .B1(n5176), .B2(n4535), .A(n5175), .ZN(n5195) );
  INV_X4 U7274 ( .A(a[4]), .ZN(n8130) );
  NAND2_X2 U7275 ( .A1(n4543), .A2(a[20]), .ZN(n6411) );
  INV_X4 U7276 ( .A(n6411), .ZN(n5178) );
  INV_X4 U7277 ( .A(a[12]), .ZN(n6553) );
  NOR2_X4 U7278 ( .A1(n5178), .A2(n5177), .ZN(n5179) );
  OAI221_X2 U7279 ( .B1(n8130), .B2(n8298), .C1(net246958), .C2(net246782), 
        .A(n5179), .ZN(n5244) );
  NAND2_X2 U7280 ( .A1(n4543), .A2(a[14]), .ZN(n7421) );
  NAND2_X2 U7281 ( .A1(net246962), .A2(a[22]), .ZN(n5181) );
  NAND2_X2 U7282 ( .A1(net247082), .A2(a[6]), .ZN(n5180) );
  NAND4_X2 U7283 ( .A1(n5314), .A2(n7421), .A3(n5181), .A4(n5180), .ZN(n5373)
         );
  AOI22_X2 U7284 ( .A1(n3977), .A2(n5244), .B1(n4561), .B2(n5373), .ZN(n5191)
         );
  NAND2_X2 U7285 ( .A1(n4543), .A2(n4578), .ZN(n7037) );
  INV_X4 U7286 ( .A(n7037), .ZN(n5183) );
  INV_X4 U7287 ( .A(a[8]), .ZN(n7240) );
  NOR2_X4 U7288 ( .A1(n5183), .A2(n5182), .ZN(n5184) );
  OAI221_X2 U7289 ( .B1(net240839), .B2(n8298), .C1(net246958), .C2(net246756), 
        .A(n5184), .ZN(n5315) );
  NAND2_X2 U7290 ( .A1(n4543), .A2(a[18]), .ZN(n6700) );
  INV_X4 U7291 ( .A(n6700), .ZN(n5186) );
  INV_X4 U7292 ( .A(a[10]), .ZN(n6901) );
  NOR2_X4 U7293 ( .A1(n5186), .A2(n5185), .ZN(n5189) );
  INV_X4 U7294 ( .A(a[2]), .ZN(n8773) );
  NAND2_X2 U7295 ( .A1(n5189), .A2(n5188), .ZN(n5273) );
  AOI22_X2 U7296 ( .A1(n4557), .A2(n5315), .B1(n4554), .B2(n5273), .ZN(n5190)
         );
  NAND2_X2 U7297 ( .A1(n5191), .A2(n5190), .ZN(n5211) );
  INV_X4 U7298 ( .A(n5211), .ZN(n5193) );
  NAND2_X2 U7299 ( .A1(net246902), .A2(a[30]), .ZN(n5236) );
  OAI22_X2 U7300 ( .A1(net245318), .A2(n5236), .B1(n620), .B2(net246782), .ZN(
        n5271) );
  NAND2_X2 U7301 ( .A1(n8318), .A2(n5271), .ZN(n5192) );
  OAI21_X4 U7302 ( .B1(n5193), .B2(n4531), .A(n5192), .ZN(n5194) );
  OAI21_X4 U7303 ( .B1(n5195), .B2(n5194), .A(n4548), .ZN(n5202) );
  NOR2_X4 U7304 ( .A1(n4551), .A2(n5196), .ZN(n5197) );
  MUX2_X2 U7305 ( .A(n4003), .B(n5197), .S(net245546), .Z(n5201) );
  NAND2_X2 U7306 ( .A1(n3988), .A2(net245541), .ZN(n5198) );
  INV_X4 U7307 ( .A(n5198), .ZN(n5666) );
  AOI221_X2 U7308 ( .B1(n5666), .B2(n8784), .C1(net247002), .C2(n3988), .A(
        n5199), .ZN(n5200) );
  NAND4_X2 U7309 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(out[28]) );
  XNOR2_X2 U7310 ( .A(n5204), .B(net246788), .ZN(n5207) );
  INV_X4 U7311 ( .A(n5205), .ZN(n5206) );
  XNOR2_X2 U7312 ( .A(n5207), .B(n5206), .ZN(n5210) );
  NOR2_X4 U7313 ( .A1(b[29]), .A2(net246788), .ZN(n5225) );
  INV_X4 U7314 ( .A(n5225), .ZN(n5208) );
  NAND2_X2 U7315 ( .A1(n5208), .A2(net245313), .ZN(n5678) );
  AOI21_X4 U7316 ( .B1(n8781), .B2(n5210), .A(n5209), .ZN(n5230) );
  INV_X4 U7317 ( .A(net245523), .ZN(net245501) );
  NAND2_X2 U7318 ( .A1(net240782), .A2(net245393), .ZN(n5229) );
  NAND2_X2 U7319 ( .A1(n4534), .A2(n5211), .ZN(n5223) );
  NAND2_X2 U7320 ( .A1(n8318), .A2(n5212), .ZN(n5222) );
  INV_X4 U7321 ( .A(n4531), .ZN(n5220) );
  NAND2_X2 U7322 ( .A1(n4558), .A2(n5787), .ZN(n5219) );
  NAND2_X2 U7323 ( .A1(n4543), .A2(a[21]), .ZN(n6283) );
  INV_X4 U7324 ( .A(n6283), .ZN(n5214) );
  INV_X4 U7325 ( .A(a[13]), .ZN(n6398) );
  NOR2_X4 U7326 ( .A1(n5214), .A2(n5213), .ZN(n5215) );
  OAI221_X2 U7327 ( .B1(n7842), .B2(n8298), .C1(net246958), .C2(net246792), 
        .A(n5215), .ZN(n5791) );
  NAND2_X2 U7328 ( .A1(n3977), .A2(n5791), .ZN(n5218) );
  NAND2_X2 U7329 ( .A1(n4555), .A2(n5788), .ZN(n5217) );
  NAND2_X2 U7330 ( .A1(n4561), .A2(n5353), .ZN(n5216) );
  NAND4_X2 U7331 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n5239)
         );
  NAND2_X2 U7332 ( .A1(n5220), .A2(n5239), .ZN(n5221) );
  NAND4_X2 U7333 ( .A1(n5224), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n5227)
         );
  NOR2_X4 U7334 ( .A1(n5225), .A2(net247049), .ZN(n5226) );
  AOI21_X4 U7335 ( .B1(n4548), .B2(n5227), .A(n5226), .ZN(n5228) );
  NAND4_X2 U7336 ( .A1(n5230), .A2(net245501), .A3(n5229), .A4(n5228), .ZN(
        out[29]) );
  INV_X4 U7337 ( .A(n5232), .ZN(n5233) );
  XNOR2_X2 U7338 ( .A(n5234), .B(n5233), .ZN(n5235) );
  NAND2_X2 U7339 ( .A1(n8781), .A2(n5235), .ZN(n5256) );
  NOR2_X4 U7340 ( .A1(n5238), .A2(n5237), .ZN(n5255) );
  INV_X4 U7341 ( .A(n5239), .ZN(n5249) );
  AOI22_X2 U7342 ( .A1(net247082), .A2(a[14]), .B1(n8834), .B2(a[6]), .ZN(
        n5242) );
  NAND2_X2 U7343 ( .A1(n4543), .A2(a[22]), .ZN(n5240) );
  INV_X4 U7344 ( .A(n5240), .ZN(n6125) );
  AOI21_X4 U7345 ( .B1(n4555), .B2(n5244), .A(n5243), .ZN(n5246) );
  AOI22_X2 U7346 ( .A1(n4561), .A2(n5315), .B1(n4557), .B2(n5273), .ZN(n5245)
         );
  NAND2_X2 U7347 ( .A1(n5246), .A2(n5245), .ZN(n5786) );
  NAND2_X2 U7348 ( .A1(n4530), .A2(n5786), .ZN(n5247) );
  OAI221_X2 U7349 ( .B1(n4535), .B2(n5249), .C1(n5248), .C2(n620), .A(n5247), 
        .ZN(n5250) );
  NAND2_X2 U7350 ( .A1(n4549), .A2(n5250), .ZN(n5254) );
  NAND2_X2 U7351 ( .A1(n3662), .A2(net245474), .ZN(n5252) );
  AOI21_X4 U7352 ( .B1(n5252), .B2(net246932), .A(n5251), .ZN(n5253) );
  NAND4_X2 U7353 ( .A1(n5256), .A2(n5255), .A3(n5254), .A4(n5253), .ZN(out[30]) );
  MUX2_X2 U7354 ( .A(n5258), .B(n5257), .S(net245465), .Z(n5263) );
  NOR2_X4 U7355 ( .A1(b[27]), .A2(net246772), .ZN(n5259) );
  INV_X4 U7356 ( .A(n5259), .ZN(n5260) );
  NAND2_X2 U7357 ( .A1(n5260), .A2(net245459), .ZN(n5682) );
  NAND2_X2 U7358 ( .A1(net247002), .A2(n5260), .ZN(n5261) );
  OAI221_X2 U7359 ( .B1(net245459), .B2(net247044), .C1(n4541), .C2(n5682), 
        .A(n5261), .ZN(n5262) );
  FA_X1 U7360 ( .A(net246772), .B(n5265), .CI(n5264), .S(n5281) );
  INV_X4 U7361 ( .A(n5267), .ZN(n5270) );
  NOR2_X4 U7362 ( .A1(net246956), .A2(n4569), .ZN(n5449) );
  NAND2_X2 U7363 ( .A1(n5449), .A2(net246908), .ZN(n5404) );
  INV_X4 U7364 ( .A(n5404), .ZN(n5268) );
  NAND2_X2 U7365 ( .A1(n5268), .A2(a[31]), .ZN(n5269) );
  AOI22_X2 U7366 ( .A1(n8318), .A2(n5301), .B1(n8841), .B2(n5271), .ZN(n5279)
         );
  NAND2_X2 U7367 ( .A1(n4554), .A2(n5315), .ZN(n5276) );
  NAND2_X2 U7368 ( .A1(n4543), .A2(a[12]), .ZN(n7827) );
  AOI21_X4 U7369 ( .B1(net247082), .B2(a[4]), .A(n5351), .ZN(n5272) );
  OAI211_X2 U7370 ( .C1(net246958), .C2(n4574), .A(n7827), .B(n5272), .ZN(
        n5424) );
  NAND2_X2 U7371 ( .A1(n4562), .A2(n5424), .ZN(n5275) );
  AOI22_X2 U7372 ( .A1(n4557), .A2(n5373), .B1(n5273), .B2(n4564), .ZN(n5274)
         );
  NAND3_X2 U7373 ( .A1(n5276), .A2(n5275), .A3(n5274), .ZN(n5302) );
  AOI22_X2 U7374 ( .A1(n8125), .A2(n5302), .B1(n8842), .B2(n5277), .ZN(n5278)
         );
  AOI21_X4 U7375 ( .B1(n4552), .B2(n5281), .A(n5280), .ZN(n5282) );
  NAND2_X2 U7376 ( .A1(n5283), .A2(n5282), .ZN(out[27]) );
  MUX2_X2 U7377 ( .A(n5286), .B(n5285), .S(n5284), .Z(n5291) );
  INV_X4 U7378 ( .A(n5287), .ZN(n5288) );
  NAND2_X2 U7379 ( .A1(n5288), .A2(net245429), .ZN(n5667) );
  NAND2_X2 U7380 ( .A1(net247002), .A2(n5288), .ZN(n5289) );
  OAI221_X2 U7381 ( .B1(net245429), .B2(net247044), .C1(n4541), .C2(n5667), 
        .A(n5289), .ZN(n5290) );
  NOR2_X4 U7382 ( .A1(n5291), .A2(n5290), .ZN(n5308) );
  FA_X1 U7383 ( .A(net246766), .B(n5293), .CI(n5292), .S(n5306) );
  AOI22_X2 U7384 ( .A1(net245389), .A2(n5295), .B1(net245348), .B2(net246908), 
        .ZN(n5323) );
  INV_X4 U7385 ( .A(n5323), .ZN(n5300) );
  NAND2_X2 U7386 ( .A1(n4543), .A2(a[11]), .ZN(n8117) );
  NAND2_X2 U7387 ( .A1(net246962), .A2(a[19]), .ZN(n5297) );
  NAND2_X2 U7388 ( .A1(net247082), .A2(a[3]), .ZN(n5296) );
  NAND4_X2 U7389 ( .A1(n5314), .A2(n8117), .A3(n5297), .A4(n5296), .ZN(n5455)
         );
  AOI22_X2 U7390 ( .A1(n5455), .A2(n4562), .B1(n4557), .B2(n5395), .ZN(n5299)
         );
  AOI22_X2 U7391 ( .A1(n4555), .A2(n5353), .B1(n5787), .B2(n4564), .ZN(n5298)
         );
  NAND2_X2 U7392 ( .A1(n5299), .A2(n5298), .ZN(n5318) );
  AOI22_X2 U7393 ( .A1(n4536), .A2(n5300), .B1(n8125), .B2(n5318), .ZN(n5304)
         );
  AOI22_X2 U7394 ( .A1(n8842), .A2(n5302), .B1(n8841), .B2(n5301), .ZN(n5303)
         );
  AOI21_X4 U7395 ( .B1(n5304), .B2(n5303), .A(n4547), .ZN(n5305) );
  AOI21_X4 U7396 ( .B1(n4552), .B2(n5306), .A(n5305), .ZN(n5307) );
  NAND2_X2 U7397 ( .A1(n5308), .A2(n5307), .ZN(out[26]) );
  XNOR2_X2 U7398 ( .A(n5311), .B(n5310), .ZN(n5329) );
  NAND2_X2 U7399 ( .A1(n4543), .A2(a[10]), .ZN(n8295) );
  NAND2_X2 U7400 ( .A1(net246962), .A2(a[18]), .ZN(n5313) );
  NAND2_X2 U7401 ( .A1(net247082), .A2(a[2]), .ZN(n5312) );
  NAND4_X2 U7402 ( .A1(n5314), .A2(n8295), .A3(n5313), .A4(n5312), .ZN(n5475)
         );
  AOI22_X2 U7403 ( .A1(n5475), .A2(n6564), .B1(n4558), .B2(n5424), .ZN(n5317)
         );
  AOI22_X2 U7404 ( .A1(n4555), .A2(n5373), .B1(n5315), .B2(n4564), .ZN(n5316)
         );
  NAND2_X2 U7405 ( .A1(n5317), .A2(n5316), .ZN(n5350) );
  AOI22_X2 U7406 ( .A1(n8125), .A2(n5350), .B1(n8842), .B2(n5318), .ZN(n5327)
         );
  INV_X4 U7407 ( .A(net245388), .ZN(net245387) );
  NAND2_X2 U7408 ( .A1(n5449), .A2(net245387), .ZN(n5320) );
  NAND2_X2 U7409 ( .A1(n5321), .A2(n5320), .ZN(n5356) );
  INV_X4 U7410 ( .A(n5356), .ZN(n5322) );
  NOR2_X4 U7411 ( .A1(n5325), .A2(n5324), .ZN(n5326) );
  AOI21_X2 U7412 ( .B1(n5327), .B2(n5326), .A(n4547), .ZN(n5328) );
  AOI21_X2 U7413 ( .B1(n4552), .B2(n5329), .A(n5328), .ZN(n5339) );
  NOR2_X4 U7414 ( .A1(n4551), .A2(n5330), .ZN(n5332) );
  MUX2_X2 U7415 ( .A(n4000), .B(n5332), .S(n5331), .Z(n5338) );
  INV_X4 U7416 ( .A(n5333), .ZN(n5335) );
  NAND2_X2 U7417 ( .A1(n5335), .A2(net245369), .ZN(n5662) );
  INV_X4 U7418 ( .A(n5662), .ZN(n5336) );
  AOI221_X2 U7419 ( .B1(n5336), .B2(n8784), .C1(net247002), .C2(n5335), .A(
        n5334), .ZN(n5337) );
  NAND3_X2 U7420 ( .A1(n5339), .A2(n5338), .A3(n5337), .ZN(out[25]) );
  MUX2_X2 U7421 ( .A(net245359), .B(n5341), .S(n4442), .Z(n5347) );
  NOR2_X4 U7422 ( .A1(b[24]), .A2(a[24]), .ZN(n5342) );
  INV_X4 U7423 ( .A(n5342), .ZN(n5343) );
  NAND2_X2 U7424 ( .A1(n5343), .A2(n5345), .ZN(n5674) );
  NAND2_X2 U7425 ( .A1(net247002), .A2(n5343), .ZN(n5344) );
  OAI221_X2 U7426 ( .B1(n5345), .B2(net247044), .C1(n4541), .C2(n5674), .A(
        n5344), .ZN(n5346) );
  NOR2_X4 U7427 ( .A1(n5347), .A2(n5346), .ZN(n5362) );
  FA_X1 U7428 ( .A(a[24]), .B(n5349), .CI(n5348), .S(n5360) );
  OAI22_X2 U7429 ( .A1(net245349), .A2(net246958), .B1(net246756), .B2(
        net245318), .ZN(n5401) );
  MUX2_X2 U7430 ( .A(n5401), .B(net245348), .S(net246902), .Z(n5380) );
  AOI22_X2 U7431 ( .A1(n8318), .A2(n5380), .B1(n8842), .B2(n5350), .ZN(n5358)
         );
  NAND2_X2 U7432 ( .A1(n4543), .A2(a[9]), .ZN(n8789) );
  AOI21_X4 U7433 ( .B1(net247082), .B2(a[1]), .A(n5351), .ZN(n5352) );
  OAI211_X2 U7434 ( .C1(net246958), .C2(n4577), .A(n8789), .B(n5352), .ZN(
        n5823) );
  AOI22_X2 U7435 ( .A1(n4561), .A2(n5823), .B1(n4558), .B2(n5455), .ZN(n5355)
         );
  AOI22_X2 U7436 ( .A1(n4555), .A2(n5395), .B1(n5353), .B2(n4564), .ZN(n5354)
         );
  NAND2_X2 U7437 ( .A1(n5355), .A2(n5354), .ZN(n5379) );
  AOI22_X2 U7438 ( .A1(n8841), .A2(n5356), .B1(n8125), .B2(n5379), .ZN(n5357)
         );
  AOI21_X4 U7439 ( .B1(n5358), .B2(n5357), .A(n4546), .ZN(n5359) );
  AOI21_X4 U7440 ( .B1(n4552), .B2(n5360), .A(n5359), .ZN(n5361) );
  NAND2_X2 U7441 ( .A1(n5362), .A2(n5361), .ZN(out[24]) );
  XNOR2_X2 U7442 ( .A(a[23]), .B(n5363), .ZN(n5364) );
  XNOR2_X2 U7443 ( .A(n5365), .B(n5364), .ZN(n5368) );
  NOR2_X4 U7444 ( .A1(b[23]), .A2(a[23]), .ZN(n5385) );
  INV_X4 U7445 ( .A(n5385), .ZN(n5366) );
  NAND2_X2 U7446 ( .A1(n5366), .A2(n6037), .ZN(n5672) );
  AOI21_X2 U7447 ( .B1(n4552), .B2(n5368), .A(n5367), .ZN(n5391) );
  NOR2_X4 U7448 ( .A1(n4551), .A2(n5369), .ZN(n5372) );
  MUX2_X2 U7449 ( .A(n5372), .B(n4004), .S(n5371), .Z(n5390) );
  AOI22_X2 U7450 ( .A1(n4561), .A2(n5474), .B1(n4558), .B2(n5475), .ZN(n5375)
         );
  AOI22_X2 U7451 ( .A1(n4555), .A2(n5424), .B1(n5373), .B2(n4564), .ZN(n5374)
         );
  NAND2_X2 U7452 ( .A1(n5375), .A2(n5374), .ZN(n5405) );
  NAND2_X2 U7453 ( .A1(n8125), .A2(n5405), .ZN(n5384) );
  NAND2_X2 U7454 ( .A1(net246962), .A2(net246902), .ZN(n5378) );
  NAND2_X2 U7455 ( .A1(n8318), .A2(n5400), .ZN(n5383) );
  NAND2_X2 U7456 ( .A1(n8842), .A2(n5379), .ZN(n5382) );
  NAND2_X2 U7457 ( .A1(n8841), .A2(n5380), .ZN(n5381) );
  NAND4_X2 U7458 ( .A1(n5384), .A2(n5383), .A3(n5382), .A4(n5381), .ZN(n5388)
         );
  AOI211_X4 U7459 ( .C1(n4548), .C2(n5388), .A(n5387), .B(n5386), .ZN(n5389)
         );
  NAND3_X2 U7460 ( .A1(n5391), .A2(n5390), .A3(n5389), .ZN(out[23]) );
  XNOR2_X2 U7461 ( .A(a[22]), .B(n5392), .ZN(n5394) );
  XNOR2_X2 U7462 ( .A(n5394), .B(n5393), .ZN(n5409) );
  NAND2_X2 U7463 ( .A1(n4558), .A2(n5823), .ZN(n5399) );
  NAND2_X2 U7464 ( .A1(n4562), .A2(n5824), .ZN(n5398) );
  NAND2_X2 U7465 ( .A1(n5395), .A2(n4565), .ZN(n5397) );
  NAND2_X2 U7466 ( .A1(n4554), .A2(n5455), .ZN(n5396) );
  NAND4_X2 U7467 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n5429)
         );
  AOI22_X2 U7468 ( .A1(n8125), .A2(n5429), .B1(n8841), .B2(n5400), .ZN(n5407)
         );
  NAND2_X2 U7469 ( .A1(n3977), .A2(n5818), .ZN(n5403) );
  NAND2_X2 U7470 ( .A1(net248516), .A2(n5401), .ZN(n5402) );
  AOI22_X2 U7471 ( .A1(n8842), .A2(n5405), .B1(n8318), .B2(n5432), .ZN(n5406)
         );
  AOI21_X2 U7472 ( .B1(n4552), .B2(n5409), .A(n5408), .ZN(n5417) );
  NOR2_X4 U7473 ( .A1(n4551), .A2(n5410), .ZN(n5412) );
  MUX2_X2 U7474 ( .A(n4001), .B(n5412), .S(n5411), .Z(n5416) );
  NAND2_X2 U7475 ( .A1(a[22]), .A2(b[22]), .ZN(n6322) );
  NAND2_X2 U7476 ( .A1(n3989), .A2(n6322), .ZN(n5589) );
  INV_X4 U7477 ( .A(n5589), .ZN(n5414) );
  AOI221_X2 U7478 ( .B1(n5414), .B2(n8784), .C1(n4267), .C2(n3989), .A(n5413), 
        .ZN(n5415) );
  NAND3_X2 U7479 ( .A1(n5417), .A2(n5416), .A3(n5415), .ZN(out[22]) );
  MUX2_X2 U7480 ( .A(net245266), .B(n5418), .S(net245268), .Z(n5421) );
  NAND2_X2 U7481 ( .A1(net246836), .A2(a[21]), .ZN(n6665) );
  NAND2_X2 U7482 ( .A1(n3993), .A2(n6665), .ZN(n5590) );
  NAND2_X2 U7483 ( .A1(n4267), .A2(n3993), .ZN(n5419) );
  OAI221_X2 U7484 ( .B1(n6665), .B2(net247044), .C1(n4541), .C2(n5590), .A(
        n5419), .ZN(n5420) );
  NOR2_X4 U7485 ( .A1(n5421), .A2(n5420), .ZN(n5438) );
  FA_X1 U7486 ( .A(a[21]), .B(n5423), .CI(n5422), .S(n5436) );
  NAND2_X2 U7487 ( .A1(n4558), .A2(n5474), .ZN(n5428) );
  NAND2_X2 U7488 ( .A1(n4562), .A2(n5994), .ZN(n5427) );
  NAND2_X2 U7489 ( .A1(n5424), .A2(n4565), .ZN(n5426) );
  NAND2_X2 U7490 ( .A1(n4554), .A2(n5475), .ZN(n5425) );
  NAND4_X2 U7491 ( .A1(n5428), .A2(n5427), .A3(n5426), .A4(n5425), .ZN(n5454)
         );
  AOI22_X2 U7492 ( .A1(n5429), .A2(n8842), .B1(n8125), .B2(n5454), .ZN(n5434)
         );
  NAND2_X2 U7493 ( .A1(n4554), .A2(n5480), .ZN(n5431) );
  INV_X4 U7494 ( .A(net245250), .ZN(net245249) );
  NAND2_X2 U7495 ( .A1(net245249), .A2(n5449), .ZN(n5430) );
  OAI211_X2 U7496 ( .C1(net248516), .C2(n5483), .A(n5431), .B(n5430), .ZN(
        n5459) );
  AOI22_X2 U7497 ( .A1(n5459), .A2(n4536), .B1(n8841), .B2(n5432), .ZN(n5433)
         );
  AOI21_X4 U7498 ( .B1(n5434), .B2(n5433), .A(n4547), .ZN(n5435) );
  AOI21_X4 U7499 ( .B1(n4552), .B2(n5436), .A(n5435), .ZN(n5437) );
  NAND2_X2 U7500 ( .A1(n5438), .A2(n5437), .ZN(out[21]) );
  MUX2_X2 U7501 ( .A(n5441), .B(n5440), .S(n4008), .Z(n5446) );
  NAND2_X2 U7502 ( .A1(a[20]), .A2(b[20]), .ZN(n6957) );
  NOR2_X4 U7503 ( .A1(a[20]), .A2(b[20]), .ZN(n5442) );
  INV_X4 U7504 ( .A(n5442), .ZN(n5443) );
  NAND2_X2 U7505 ( .A1(n5443), .A2(n6957), .ZN(n5593) );
  NAND2_X2 U7506 ( .A1(n4267), .A2(n5443), .ZN(n5444) );
  OAI221_X2 U7507 ( .B1(n6957), .B2(net247044), .C1(n4541), .C2(n5593), .A(
        n5444), .ZN(n5445) );
  FA_X1 U7508 ( .A(a[20]), .B(n5448), .CI(n5447), .S(n5463) );
  INV_X4 U7509 ( .A(n5449), .ZN(n5453) );
  AOI22_X2 U7510 ( .A1(n5450), .A2(n4569), .B1(n5449), .B2(a[24]), .ZN(n5821)
         );
  NAND2_X2 U7511 ( .A1(n4554), .A2(n5818), .ZN(n5451) );
  AOI22_X2 U7512 ( .A1(n5454), .A2(n8842), .B1(n8318), .B2(n5484), .ZN(n5461)
         );
  NAND2_X2 U7513 ( .A1(n5455), .A2(n4565), .ZN(n5458) );
  NAND2_X2 U7514 ( .A1(n4554), .A2(n5823), .ZN(n5457) );
  AOI22_X2 U7515 ( .A1(n4561), .A2(n6129), .B1(n4557), .B2(n5824), .ZN(n5456)
         );
  NAND3_X2 U7516 ( .A1(n5458), .A2(n5457), .A3(n5456), .ZN(n5485) );
  AOI22_X2 U7517 ( .A1(n8125), .A2(n5485), .B1(n8841), .B2(n5459), .ZN(n5460)
         );
  NAND2_X2 U7518 ( .A1(n5465), .A2(n5464), .ZN(out[20]) );
  MUX2_X2 U7519 ( .A(net245207), .B(n5466), .S(net245209), .Z(n5471) );
  NAND2_X2 U7520 ( .A1(b[19]), .A2(a[19]), .ZN(n7458) );
  NOR2_X4 U7521 ( .A1(a[19]), .A2(b[19]), .ZN(n5467) );
  INV_X4 U7522 ( .A(n5467), .ZN(n5468) );
  NAND2_X2 U7523 ( .A1(n5468), .A2(n7458), .ZN(n5575) );
  NAND2_X2 U7524 ( .A1(n4267), .A2(n5468), .ZN(n5469) );
  OAI221_X2 U7525 ( .B1(n7458), .B2(net247044), .C1(n4541), .C2(n5575), .A(
        n5469), .ZN(n5470) );
  NOR2_X4 U7526 ( .A1(n5471), .A2(n5470), .ZN(n5491) );
  FA_X1 U7527 ( .A(a[19]), .B(n5473), .CI(n5472), .S(n5489) );
  NAND2_X2 U7528 ( .A1(n4554), .A2(n5474), .ZN(n5479) );
  NAND2_X2 U7529 ( .A1(n4558), .A2(n5994), .ZN(n5478) );
  NAND2_X2 U7530 ( .A1(n5475), .A2(n4565), .ZN(n5477) );
  NAND2_X2 U7531 ( .A1(n4562), .A2(n6273), .ZN(n5476) );
  NAND4_X2 U7532 ( .A1(n5479), .A2(n5478), .A3(n5477), .A4(n5476), .ZN(n5828)
         );
  NAND2_X2 U7533 ( .A1(n4558), .A2(n5480), .ZN(n5482) );
  NAND2_X2 U7534 ( .A1(n6280), .A2(n4565), .ZN(n5481) );
  OAI211_X2 U7535 ( .C1(n5483), .C2(net246908), .A(n5482), .B(n5481), .ZN(
        n5822) );
  AOI22_X2 U7536 ( .A1(n8125), .A2(n5828), .B1(n8318), .B2(n5822), .ZN(n5487)
         );
  AOI22_X2 U7537 ( .A1(n8842), .A2(n5485), .B1(n8841), .B2(n5484), .ZN(n5486)
         );
  AOI21_X4 U7538 ( .B1(n5487), .B2(n5486), .A(n4547), .ZN(n5488) );
  AOI21_X4 U7539 ( .B1(n4552), .B2(n5489), .A(n5488), .ZN(n5490) );
  NAND2_X2 U7540 ( .A1(n5491), .A2(n5490), .ZN(out[19]) );
  INV_X4 U7541 ( .A(n5748), .ZN(n5661) );
  NAND2_X2 U7542 ( .A1(b[3]), .A2(n8289), .ZN(n5732) );
  NAND2_X2 U7543 ( .A1(a[3]), .A2(n8281), .ZN(n5625) );
  NAND2_X2 U7544 ( .A1(n5732), .A2(n5625), .ZN(n8137) );
  INV_X4 U7545 ( .A(n8137), .ZN(n5747) );
  XNOR2_X2 U7546 ( .A(a[2]), .B(b[2]), .ZN(n5733) );
  NAND2_X2 U7547 ( .A1(n5747), .A2(n5733), .ZN(n5538) );
  NAND2_X2 U7548 ( .A1(n5733), .A2(n5625), .ZN(n5492) );
  NAND2_X2 U7549 ( .A1(n5492), .A2(n8137), .ZN(n5537) );
  NAND2_X2 U7550 ( .A1(a[7]), .A2(net242655), .ZN(n5618) );
  INV_X4 U7551 ( .A(n5618), .ZN(n5535) );
  NAND2_X2 U7552 ( .A1(b[10]), .A2(n6901), .ZN(n5609) );
  INV_X4 U7553 ( .A(b[14]), .ZN(net244239) );
  NOR2_X4 U7554 ( .A1(b[15]), .A2(n4580), .ZN(n5527) );
  NOR2_X4 U7555 ( .A1(b[17]), .A2(n4577), .ZN(n5523) );
  INV_X4 U7556 ( .A(b[18]), .ZN(net244808) );
  NOR2_X4 U7557 ( .A1(a[18]), .A2(net244808), .ZN(n5521) );
  NOR2_X4 U7558 ( .A1(b[19]), .A2(n4575), .ZN(n5519) );
  NOR2_X4 U7559 ( .A1(a[20]), .A2(net246832), .ZN(n5517) );
  NOR2_X4 U7560 ( .A1(a[23]), .A2(net246850), .ZN(n5510) );
  NOR2_X4 U7561 ( .A1(net248516), .A2(net246804), .ZN(n5494) );
  NAND2_X2 U7562 ( .A1(net249231), .A2(net246812), .ZN(n5680) );
  NAND2_X2 U7563 ( .A1(net248517), .A2(net246804), .ZN(n5493) );
  OAI21_X4 U7564 ( .B1(n5494), .B2(n5680), .A(n5493), .ZN(n5679) );
  NAND2_X2 U7565 ( .A1(net246788), .A2(n4569), .ZN(n5495) );
  OAI21_X4 U7566 ( .B1(n5496), .B2(n5679), .A(n5495), .ZN(n5664) );
  NAND2_X2 U7567 ( .A1(net246878), .A2(net246782), .ZN(n5497) );
  OAI21_X4 U7568 ( .B1(n5498), .B2(n5664), .A(n5497), .ZN(n5683) );
  NAND2_X2 U7569 ( .A1(net246772), .A2(net246874), .ZN(n5499) );
  OAI21_X4 U7570 ( .B1(n5500), .B2(n5683), .A(n5499), .ZN(n5501) );
  INV_X4 U7571 ( .A(n5501), .ZN(n5668) );
  NAND2_X2 U7572 ( .A1(net246766), .A2(net246868), .ZN(n5502) );
  OAI21_X4 U7573 ( .B1(n5668), .B2(n5503), .A(n5502), .ZN(n5663) );
  OAI21_X4 U7574 ( .B1(n5505), .B2(n5663), .A(n5504), .ZN(n5675) );
  INV_X4 U7575 ( .A(n5675), .ZN(n5508) );
  NOR2_X4 U7576 ( .A1(b[24]), .A2(net246756), .ZN(n5507) );
  NAND2_X2 U7577 ( .A1(b[24]), .A2(net246756), .ZN(n5506) );
  OAI21_X4 U7578 ( .B1(n5508), .B2(n5507), .A(n5506), .ZN(n5673) );
  NAND2_X2 U7579 ( .A1(a[23]), .A2(net246850), .ZN(n5509) );
  OAI21_X4 U7580 ( .B1(n5510), .B2(n5673), .A(n5509), .ZN(n5588) );
  INV_X4 U7581 ( .A(n5588), .ZN(n5513) );
  NOR2_X4 U7582 ( .A1(a[22]), .A2(net246844), .ZN(n5512) );
  NAND2_X2 U7583 ( .A1(a[22]), .A2(net246844), .ZN(n5511) );
  OAI21_X4 U7584 ( .B1(n5513), .B2(n5512), .A(n5511), .ZN(n5591) );
  NAND2_X2 U7585 ( .A1(net246836), .A2(n4572), .ZN(n5514) );
  OAI21_X4 U7586 ( .B1(n5515), .B2(n5591), .A(n5514), .ZN(n5594) );
  NAND2_X2 U7587 ( .A1(a[20]), .A2(net246832), .ZN(n5516) );
  OAI21_X4 U7588 ( .B1(n5517), .B2(n5594), .A(n5516), .ZN(n5576) );
  NAND2_X2 U7589 ( .A1(b[19]), .A2(n4575), .ZN(n5518) );
  OAI21_X4 U7590 ( .B1(n5519), .B2(n5576), .A(n5518), .ZN(n5592) );
  NAND2_X2 U7591 ( .A1(a[18]), .A2(net244808), .ZN(n5520) );
  OAI21_X4 U7592 ( .B1(n5521), .B2(n5592), .A(n5520), .ZN(n5574) );
  NAND2_X2 U7593 ( .A1(b[17]), .A2(n4577), .ZN(n5522) );
  OAI21_X4 U7594 ( .B1(n5523), .B2(n5574), .A(n5522), .ZN(n5572) );
  NAND2_X2 U7595 ( .A1(a[16]), .A2(net244627), .ZN(n5524) );
  OAI21_X4 U7596 ( .B1(n5525), .B2(n5572), .A(n5524), .ZN(n5564) );
  NAND2_X2 U7597 ( .A1(b[15]), .A2(n4580), .ZN(n5526) );
  OAI21_X4 U7598 ( .B1(n5527), .B2(n5564), .A(n5526), .ZN(n5562) );
  NAND2_X2 U7599 ( .A1(a[14]), .A2(net244239), .ZN(n5528) );
  OAI21_X4 U7600 ( .B1(n5529), .B2(n5562), .A(n5528), .ZN(n5563) );
  INV_X4 U7601 ( .A(n5563), .ZN(n5531) );
  INV_X4 U7602 ( .A(b[13]), .ZN(n6389) );
  NAND2_X2 U7603 ( .A1(a[13]), .A2(n6389), .ZN(n5530) );
  AOI22_X2 U7604 ( .A1(n5531), .A2(n5530), .B1(b[13]), .B2(n6398), .ZN(n5565)
         );
  NAND2_X2 U7605 ( .A1(b[12]), .A2(n6553), .ZN(n5532) );
  INV_X4 U7606 ( .A(b[12]), .ZN(net243844) );
  AOI22_X2 U7607 ( .A1(n5565), .A2(n5532), .B1(a[12]), .B2(net243844), .ZN(
        n5587) );
  INV_X4 U7608 ( .A(b[11]), .ZN(net243628) );
  NAND2_X2 U7609 ( .A1(a[11]), .A2(net243628), .ZN(n5585) );
  NAND2_X2 U7610 ( .A1(n5587), .A2(n5585), .ZN(n5611) );
  INV_X4 U7611 ( .A(b[10]), .ZN(net243587) );
  NAND2_X2 U7612 ( .A1(a[10]), .A2(net243587), .ZN(n5612) );
  INV_X4 U7613 ( .A(n5612), .ZN(n5533) );
  AOI21_X4 U7614 ( .B1(n5609), .B2(n5611), .A(n5533), .ZN(n5551) );
  INV_X4 U7615 ( .A(b[9]), .ZN(net243356) );
  NAND2_X2 U7616 ( .A1(a[9]), .A2(net243356), .ZN(n5614) );
  NAND2_X2 U7617 ( .A1(a[8]), .A2(net242878), .ZN(n5616) );
  INV_X4 U7618 ( .A(b[6]), .ZN(n7404) );
  NAND2_X2 U7619 ( .A1(a[6]), .A2(n7404), .ZN(n5619) );
  INV_X4 U7620 ( .A(n5619), .ZN(n5534) );
  NOR3_X4 U7621 ( .A1(n5535), .A2(n5555), .A3(n5534), .ZN(n5546) );
  INV_X4 U7622 ( .A(b[4]), .ZN(net242110) );
  NAND2_X2 U7623 ( .A1(a[4]), .A2(net242110), .ZN(n5623) );
  INV_X4 U7624 ( .A(b[5]), .ZN(net242361) );
  NAND2_X2 U7625 ( .A1(a[5]), .A2(net242361), .ZN(n5621) );
  INV_X4 U7626 ( .A(n5539), .ZN(n5536) );
  MUX2_X2 U7627 ( .A(n5538), .B(n5537), .S(n5536), .Z(n5545) );
  NAND2_X2 U7628 ( .A1(b[1]), .A2(net240852), .ZN(n5734) );
  NAND2_X2 U7629 ( .A1(n5734), .A2(net245029), .ZN(n8783) );
  INV_X4 U7630 ( .A(n8783), .ZN(n5745) );
  NAND2_X2 U7631 ( .A1(b[0]), .A2(net240839), .ZN(n5776) );
  NAND2_X2 U7632 ( .A1(n5776), .A2(net244873), .ZN(n5629) );
  INV_X4 U7633 ( .A(n5629), .ZN(n8851) );
  NAND2_X2 U7634 ( .A1(n5745), .A2(n8851), .ZN(n5543) );
  NAND2_X2 U7635 ( .A1(n8851), .A2(net245029), .ZN(n5736) );
  NAND2_X2 U7636 ( .A1(n5736), .A2(n8783), .ZN(n5542) );
  INV_X4 U7637 ( .A(b[2]), .ZN(net241554) );
  NAND2_X2 U7638 ( .A1(a[2]), .A2(net241554), .ZN(n5626) );
  INV_X4 U7639 ( .A(n5626), .ZN(n5540) );
  INV_X4 U7640 ( .A(n5625), .ZN(n5582) );
  NOR3_X4 U7641 ( .A1(n5540), .A2(n5582), .A3(n5539), .ZN(n5541) );
  MUX2_X2 U7642 ( .A(n5543), .B(n5542), .S(n5541), .Z(n5544) );
  NAND2_X2 U7643 ( .A1(b[5]), .A2(n7842), .ZN(n5737) );
  NAND2_X2 U7644 ( .A1(n5737), .A2(n5621), .ZN(n7647) );
  INV_X4 U7645 ( .A(n7647), .ZN(n5760) );
  NAND2_X2 U7646 ( .A1(b[4]), .A2(n8130), .ZN(n5746) );
  NAND2_X2 U7647 ( .A1(n5746), .A2(n5623), .ZN(n7848) );
  INV_X4 U7648 ( .A(n7848), .ZN(n5740) );
  NAND2_X2 U7649 ( .A1(n5760), .A2(n5740), .ZN(n5548) );
  NAND2_X2 U7650 ( .A1(n5740), .A2(n5621), .ZN(n5739) );
  NAND2_X2 U7651 ( .A1(n5739), .A2(n7647), .ZN(n5547) );
  MUX2_X2 U7652 ( .A(n5548), .B(n5547), .S(n5546), .Z(n5561) );
  NAND2_X2 U7653 ( .A1(b[9]), .A2(n7029), .ZN(n5727) );
  NAND2_X2 U7654 ( .A1(n5727), .A2(n5614), .ZN(n6900) );
  INV_X4 U7655 ( .A(n6900), .ZN(n5549) );
  XNOR2_X2 U7656 ( .A(a[8]), .B(b[8]), .ZN(n5728) );
  NAND2_X2 U7657 ( .A1(n5549), .A2(n5728), .ZN(n5553) );
  NAND2_X2 U7658 ( .A1(n5728), .A2(n5614), .ZN(n5550) );
  NAND2_X2 U7659 ( .A1(n5550), .A2(n6900), .ZN(n5552) );
  MUX2_X2 U7660 ( .A(n5553), .B(n5552), .S(n5551), .Z(n5560) );
  INV_X4 U7661 ( .A(a[7]), .ZN(n7409) );
  NAND2_X2 U7662 ( .A1(b[7]), .A2(n7409), .ZN(n5724) );
  NAND2_X2 U7663 ( .A1(n5724), .A2(n5618), .ZN(n7239) );
  INV_X4 U7664 ( .A(n7239), .ZN(n5554) );
  INV_X4 U7665 ( .A(a[6]), .ZN(n7648) );
  NAND2_X2 U7666 ( .A1(b[6]), .A2(n7648), .ZN(n5759) );
  NAND2_X2 U7667 ( .A1(n5759), .A2(n5619), .ZN(n7407) );
  INV_X4 U7668 ( .A(n7407), .ZN(n5644) );
  NAND2_X2 U7669 ( .A1(n5554), .A2(n5644), .ZN(n5558) );
  NAND2_X2 U7670 ( .A1(n5644), .A2(n5618), .ZN(n5723) );
  NAND2_X2 U7671 ( .A1(n5723), .A2(n7239), .ZN(n5557) );
  INV_X4 U7672 ( .A(n5555), .ZN(n5556) );
  MUX2_X2 U7673 ( .A(n5558), .B(n5557), .S(n5556), .Z(n5559) );
  XNOR2_X2 U7674 ( .A(a[14]), .B(b[14]), .ZN(n6114) );
  XNOR2_X2 U7675 ( .A(n5562), .B(n6114), .ZN(n5570) );
  XNOR2_X2 U7676 ( .A(b[13]), .B(a[13]), .ZN(n6262) );
  XNOR2_X2 U7677 ( .A(n6262), .B(n5563), .ZN(n5568) );
  XNOR2_X2 U7678 ( .A(b[15]), .B(a[15]), .ZN(n5973) );
  XNOR2_X2 U7679 ( .A(n5564), .B(n5973), .ZN(n5567) );
  XNOR2_X2 U7680 ( .A(b[12]), .B(a[12]), .ZN(n6395) );
  XNOR2_X2 U7681 ( .A(n5565), .B(n6395), .ZN(n5566) );
  NOR2_X4 U7682 ( .A1(n5570), .A2(n5569), .ZN(n5651) );
  XOR2_X2 U7683 ( .A(n5572), .B(n5571), .Z(n5579) );
  NOR2_X4 U7684 ( .A1(b[17]), .A2(a[17]), .ZN(n5573) );
  INV_X4 U7685 ( .A(n5573), .ZN(n5859) );
  NAND2_X2 U7686 ( .A1(b[17]), .A2(a[17]), .ZN(n8182) );
  NAND2_X2 U7687 ( .A1(n5859), .A2(n8182), .ZN(n5857) );
  XNOR2_X2 U7688 ( .A(n5574), .B(n5857), .ZN(n5578) );
  XNOR2_X2 U7689 ( .A(n5576), .B(n5575), .ZN(n5577) );
  INV_X4 U7690 ( .A(n5649), .ZN(n5580) );
  NAND2_X2 U7691 ( .A1(n5651), .A2(n5580), .ZN(n5581) );
  INV_X4 U7692 ( .A(n5581), .ZN(n5768) );
  INV_X4 U7693 ( .A(n5733), .ZN(n8287) );
  NAND2_X2 U7694 ( .A1(n5582), .A2(n8287), .ZN(n5583) );
  OAI221_X2 U7695 ( .B1(n8851), .B2(net245029), .C1(n5740), .C2(n5621), .A(
        n5583), .ZN(n5766) );
  INV_X4 U7696 ( .A(n5766), .ZN(n5584) );
  NAND2_X2 U7697 ( .A1(n5768), .A2(n5584), .ZN(n5605) );
  NAND2_X2 U7698 ( .A1(n5609), .A2(n5612), .ZN(n6718) );
  XNOR2_X2 U7699 ( .A(n6718), .B(n5611), .ZN(n5604) );
  INV_X4 U7700 ( .A(n5728), .ZN(n7027) );
  NAND2_X2 U7701 ( .A1(n5615), .A2(n7027), .ZN(n5603) );
  NAND2_X2 U7702 ( .A1(b[11]), .A2(n6712), .ZN(n5610) );
  NAND2_X2 U7703 ( .A1(n5585), .A2(n5610), .ZN(n6552) );
  INV_X4 U7704 ( .A(n6552), .ZN(n5586) );
  XNOR2_X2 U7705 ( .A(n5587), .B(n5586), .ZN(n5694) );
  INV_X4 U7706 ( .A(n5694), .ZN(n5602) );
  NAND2_X2 U7707 ( .A1(n5535), .A2(n7407), .ZN(n5601) );
  XNOR2_X2 U7708 ( .A(n5589), .B(n5588), .ZN(n5599) );
  XNOR2_X2 U7709 ( .A(n5591), .B(n5590), .ZN(n5598) );
  NAND2_X2 U7710 ( .A1(a[18]), .A2(b[18]), .ZN(n7767) );
  NAND2_X2 U7711 ( .A1(n3990), .A2(n7767), .ZN(n5837) );
  XOR2_X2 U7712 ( .A(n5592), .B(n5837), .Z(n5597) );
  INV_X4 U7713 ( .A(n5593), .ZN(n5595) );
  XNOR2_X2 U7714 ( .A(n5595), .B(n5594), .ZN(n5596) );
  NAND4_X2 U7715 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n5697)
         );
  INV_X4 U7716 ( .A(n5697), .ZN(n5600) );
  NAND4_X2 U7717 ( .A1(n5603), .A2(n5602), .A3(n5601), .A4(n5600), .ZN(n5769)
         );
  NAND4_X2 U7718 ( .A1(n5608), .A2(net245052), .A3(n5607), .A4(n5606), .ZN(
        n5659) );
  INV_X4 U7719 ( .A(n5746), .ZN(n5624) );
  INV_X4 U7720 ( .A(n5759), .ZN(n5620) );
  INV_X4 U7721 ( .A(n5609), .ZN(n5613) );
  NAND2_X2 U7722 ( .A1(n5611), .A2(n5610), .ZN(n5630) );
  OAI21_X4 U7723 ( .B1(n5613), .B2(n5630), .A(n5612), .ZN(n5638) );
  INV_X4 U7724 ( .A(n5614), .ZN(n5615) );
  AOI21_X4 U7725 ( .B1(n5638), .B2(n5727), .A(n5615), .ZN(n5633) );
  NAND2_X2 U7726 ( .A1(b[8]), .A2(n7240), .ZN(n5756) );
  INV_X4 U7727 ( .A(n5756), .ZN(n5617) );
  OAI21_X4 U7728 ( .B1(n5633), .B2(n5617), .A(n5616), .ZN(n5646) );
  AOI21_X4 U7729 ( .B1(n5646), .B2(n5724), .A(n5535), .ZN(n5645) );
  OAI21_X4 U7730 ( .B1(n5620), .B2(n5645), .A(n5619), .ZN(n5643) );
  INV_X4 U7731 ( .A(n5621), .ZN(n5622) );
  AOI21_X4 U7732 ( .B1(n5643), .B2(n5737), .A(n5622), .ZN(n5637) );
  OAI21_X4 U7733 ( .B1(n5624), .B2(n5637), .A(n5623), .ZN(n5641) );
  AOI21_X4 U7734 ( .B1(n5641), .B2(n5732), .A(n5582), .ZN(n5634) );
  NAND2_X2 U7735 ( .A1(b[2]), .A2(n8773), .ZN(n5744) );
  INV_X4 U7736 ( .A(n5744), .ZN(n5627) );
  OAI21_X4 U7737 ( .B1(n5634), .B2(n5627), .A(n5626), .ZN(n5642) );
  NAND2_X2 U7738 ( .A1(n5642), .A2(n5734), .ZN(n5628) );
  NAND2_X2 U7739 ( .A1(n5628), .A2(net245029), .ZN(n5777) );
  NAND2_X2 U7740 ( .A1(n5777), .A2(n5629), .ZN(n5706) );
  INV_X4 U7741 ( .A(n5706), .ZN(n5632) );
  XNOR2_X2 U7742 ( .A(n6718), .B(n5630), .ZN(n5754) );
  INV_X4 U7743 ( .A(n5754), .ZN(n5631) );
  XNOR2_X2 U7744 ( .A(n5633), .B(n7027), .ZN(n5707) );
  INV_X4 U7745 ( .A(n5707), .ZN(n5636) );
  XNOR2_X2 U7746 ( .A(n5634), .B(n8287), .ZN(n5705) );
  INV_X4 U7747 ( .A(n5705), .ZN(n5635) );
  XNOR2_X2 U7748 ( .A(n5637), .B(n7848), .ZN(n5640) );
  XNOR2_X2 U7749 ( .A(n6900), .B(n5638), .ZN(n5758) );
  INV_X4 U7750 ( .A(n5758), .ZN(n5639) );
  NAND2_X2 U7751 ( .A1(n5640), .A2(n5639), .ZN(n5709) );
  XNOR2_X2 U7752 ( .A(n8137), .B(n5641), .ZN(n5710) );
  XNOR2_X2 U7753 ( .A(n5642), .B(n8783), .ZN(n5708) );
  XNOR2_X2 U7754 ( .A(n5645), .B(n5644), .ZN(n5691) );
  INV_X4 U7755 ( .A(n5691), .ZN(n5648) );
  XNOR2_X2 U7756 ( .A(n7239), .B(n5646), .ZN(n5692) );
  NAND3_X2 U7757 ( .A1(n3905), .A2(n5648), .A3(n5647), .ZN(n5653) );
  NAND3_X2 U7758 ( .A1(n5651), .A2(ALUCtrl[2]), .A3(n5650), .ZN(n5652) );
  NAND4_X2 U7759 ( .A1(n5657), .A2(n5656), .A3(n5655), .A4(n5654), .ZN(n5658)
         );
  MUX2_X2 U7760 ( .A(n5659), .B(n5658), .S(ALUCtrl[3]), .Z(n5660) );
  XNOR2_X2 U7761 ( .A(n5663), .B(n5662), .ZN(n5703) );
  INV_X4 U7762 ( .A(n5664), .ZN(n5665) );
  XNOR2_X2 U7763 ( .A(n5666), .B(n5665), .ZN(n5704) );
  INV_X4 U7764 ( .A(n5704), .ZN(n5671) );
  INV_X4 U7765 ( .A(n5667), .ZN(n5669) );
  XNOR2_X2 U7766 ( .A(n5669), .B(n5668), .ZN(n5702) );
  INV_X4 U7767 ( .A(n5702), .ZN(n5670) );
  XNOR2_X2 U7768 ( .A(n5673), .B(n5672), .ZN(n5764) );
  INV_X4 U7769 ( .A(n5764), .ZN(n5677) );
  XNOR2_X2 U7770 ( .A(n5675), .B(n5674), .ZN(n5676) );
  INV_X4 U7771 ( .A(n5676), .ZN(n5762) );
  NAND2_X2 U7772 ( .A1(n5677), .A2(n5762), .ZN(n5693) );
  XNOR2_X2 U7773 ( .A(n5679), .B(n5678), .ZN(n5770) );
  NAND2_X2 U7774 ( .A1(a[31]), .A2(net246918), .ZN(n5681) );
  NAND2_X2 U7775 ( .A1(n5681), .A2(n5680), .ZN(n5765) );
  INV_X4 U7776 ( .A(n5682), .ZN(n5685) );
  INV_X4 U7777 ( .A(n5683), .ZN(n5684) );
  XNOR2_X2 U7778 ( .A(n5685), .B(n5684), .ZN(n5698) );
  INV_X4 U7779 ( .A(n5698), .ZN(n5761) );
  NAND2_X2 U7780 ( .A1(n5686), .A2(n5761), .ZN(n5687) );
  NAND4_X2 U7781 ( .A1(n5690), .A2(n5703), .A3(n5689), .A4(n5688), .ZN(n5722)
         );
  NOR2_X4 U7782 ( .A1(n5692), .A2(n5691), .ZN(n5696) );
  INV_X4 U7783 ( .A(n5765), .ZN(n5808) );
  NAND3_X2 U7784 ( .A1(n5768), .A2(n5808), .A3(n5699), .ZN(n5700) );
  NOR2_X4 U7785 ( .A1(n5701), .A2(n5700), .ZN(n5716) );
  NAND4_X2 U7786 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n3985), .ZN(n5714)
         );
  INV_X4 U7787 ( .A(n5708), .ZN(n5712) );
  NOR2_X4 U7788 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  NAND4_X2 U7789 ( .A1(n5712), .A2(n5748), .A3(n5754), .A4(n5711), .ZN(n5713)
         );
  NOR2_X4 U7790 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  INV_X4 U7791 ( .A(n5777), .ZN(n5718) );
  INV_X4 U7792 ( .A(n5776), .ZN(n5717) );
  AOI21_X4 U7793 ( .B1(n5718), .B2(net244873), .A(n5717), .ZN(n5780) );
  MUX2_X2 U7794 ( .A(ALUCtrl[2]), .B(n5719), .S(n5780), .Z(n5720) );
  NAND2_X2 U7795 ( .A1(n5720), .A2(net244933), .ZN(n5721) );
  MUX2_X2 U7796 ( .A(n5722), .B(n5721), .S(ALUCtrl[1]), .Z(n5784) );
  INV_X4 U7797 ( .A(n5723), .ZN(n5726) );
  INV_X4 U7798 ( .A(n5724), .ZN(n5725) );
  MUX2_X2 U7799 ( .A(n7407), .B(n5726), .S(n5725), .Z(n5731) );
  INV_X4 U7800 ( .A(n5727), .ZN(n5729) );
  XNOR2_X2 U7801 ( .A(n5729), .B(n5728), .ZN(n5730) );
  NOR2_X4 U7802 ( .A1(n5731), .A2(n5730), .ZN(n5755) );
  XNOR2_X2 U7803 ( .A(n5733), .B(n5732), .ZN(n5743) );
  INV_X4 U7804 ( .A(n5734), .ZN(n5735) );
  MUX2_X2 U7805 ( .A(n8851), .B(n5736), .S(n5735), .Z(n5742) );
  INV_X4 U7806 ( .A(n5737), .ZN(n5738) );
  MUX2_X2 U7807 ( .A(n5740), .B(n5739), .S(n5738), .Z(n5741) );
  NAND3_X2 U7808 ( .A1(n5743), .A2(n5742), .A3(n5741), .ZN(n5752) );
  XNOR2_X2 U7809 ( .A(n5745), .B(n5744), .ZN(n5750) );
  XNOR2_X2 U7810 ( .A(n5747), .B(n5746), .ZN(n5749) );
  NAND3_X2 U7811 ( .A1(n5750), .A2(n5749), .A3(n5748), .ZN(n5751) );
  NOR2_X4 U7812 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  NAND4_X2 U7813 ( .A1(n5755), .A2(n5754), .A3(n3985), .A4(n5753), .ZN(
        net244874) );
  XNOR2_X2 U7814 ( .A(n7239), .B(n5756), .ZN(n5757) );
  NOR2_X4 U7815 ( .A1(n5758), .A2(n5757), .ZN(n5775) );
  XNOR2_X2 U7816 ( .A(n5760), .B(n5759), .ZN(n5774) );
  NAND2_X2 U7817 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  NOR2_X4 U7818 ( .A1(n5764), .A2(n5763), .ZN(n5773) );
  NAND2_X2 U7819 ( .A1(n5768), .A2(n5767), .ZN(n5771) );
  NAND4_X2 U7820 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .ZN(
        net244875) );
  INV_X4 U7821 ( .A(net244873), .ZN(net244872) );
  AOI21_X2 U7822 ( .B1(n5777), .B2(n5776), .A(net244872), .ZN(n5779) );
  NOR2_X4 U7823 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  NAND3_X2 U7824 ( .A1(n5784), .A2(net244862), .A3(n5783), .ZN(n5785) );
  INV_X4 U7825 ( .A(n5785), .ZN(n5814) );
  INV_X4 U7826 ( .A(n5786), .ZN(n5800) );
  INV_X4 U7827 ( .A(n5787), .ZN(n5790) );
  NAND2_X2 U7828 ( .A1(n4558), .A2(n5788), .ZN(n5789) );
  INV_X4 U7829 ( .A(n5791), .ZN(n5796) );
  NAND2_X2 U7830 ( .A1(n8834), .A2(a[7]), .ZN(n5793) );
  NAND2_X2 U7831 ( .A1(net247082), .A2(a[15]), .ZN(n5792) );
  NAND2_X2 U7832 ( .A1(n4543), .A2(a[23]), .ZN(n5986) );
  NAND3_X2 U7833 ( .A1(n5793), .A2(n5792), .A3(n5986), .ZN(n5794) );
  NAND2_X2 U7834 ( .A1(n5794), .A2(n4565), .ZN(n5795) );
  AOI21_X4 U7835 ( .B1(n4548), .B2(n5802), .A(n5801), .ZN(n5813) );
  NAND3_X2 U7836 ( .A1(n1671), .A2(n4549), .A3(net246918), .ZN(n5804) );
  NAND3_X2 U7837 ( .A1(n8841), .A2(net244841), .A3(net246932), .ZN(n5803) );
  NAND3_X2 U7838 ( .A1(n5804), .A2(net247048), .A3(n5803), .ZN(n5811) );
  XNOR2_X2 U7839 ( .A(net246926), .B(a[31]), .ZN(n5806) );
  XNOR2_X2 U7840 ( .A(n5806), .B(n5805), .ZN(n5807) );
  NOR2_X2 U7841 ( .A1(n5807), .A2(n8856), .ZN(n5810) );
  AOI211_X4 U7842 ( .C1(a[31]), .C2(n5811), .A(n5810), .B(n5809), .ZN(n5812)
         );
  OAI211_X2 U7843 ( .C1(n5814), .C2(net246932), .A(n5813), .B(n5812), .ZN(
        out[31]) );
  XNOR2_X2 U7844 ( .A(a[18]), .B(n5815), .ZN(n5817) );
  XNOR2_X2 U7845 ( .A(n5817), .B(n5816), .ZN(n5832) );
  NAND2_X2 U7846 ( .A1(n4558), .A2(n5818), .ZN(n5820) );
  NAND2_X2 U7847 ( .A1(n6408), .A2(n4565), .ZN(n5819) );
  OAI211_X2 U7848 ( .C1(n5821), .C2(net246908), .A(n5820), .B(n5819), .ZN(
        n5847) );
  AOI22_X2 U7849 ( .A1(n8841), .A2(n5822), .B1(n8318), .B2(n5847), .ZN(n5830)
         );
  NAND2_X2 U7850 ( .A1(n5823), .A2(n4565), .ZN(n5827) );
  NAND2_X2 U7851 ( .A1(n4562), .A2(n6404), .ZN(n5826) );
  AOI22_X2 U7852 ( .A1(n4557), .A2(n6129), .B1(n4555), .B2(n5824), .ZN(n5825)
         );
  NAND3_X2 U7853 ( .A1(n5827), .A2(n5826), .A3(n5825), .ZN(n5846) );
  AOI22_X2 U7854 ( .A1(n8125), .A2(n5846), .B1(n8842), .B2(n5828), .ZN(n5829)
         );
  AOI21_X2 U7855 ( .B1(n5830), .B2(n5829), .A(n4547), .ZN(n5831) );
  AOI21_X2 U7856 ( .B1(n4552), .B2(n5832), .A(n5831), .ZN(n5842) );
  NOR2_X4 U7857 ( .A1(n4551), .A2(n5833), .ZN(n5836) );
  MUX2_X2 U7858 ( .A(n5836), .B(n4005), .S(n5835), .Z(n5841) );
  INV_X4 U7859 ( .A(n5837), .ZN(n5839) );
  AOI221_X2 U7860 ( .B1(n5839), .B2(n8784), .C1(n4267), .C2(n3990), .A(n5838), 
        .ZN(n5840) );
  NAND3_X2 U7861 ( .A1(n5842), .A2(n5841), .A3(n5840), .ZN(out[18]) );
  XNOR2_X2 U7862 ( .A(a[17]), .B(n5843), .ZN(n5844) );
  XNOR2_X2 U7863 ( .A(n5845), .B(n5844), .ZN(n5853) );
  AOI22_X2 U7864 ( .A1(n8841), .A2(n5847), .B1(n8842), .B2(n5846), .ZN(n5851)
         );
  AOI22_X2 U7865 ( .A1(n8125), .A2(n5849), .B1(n8318), .B2(n5848), .ZN(n5850)
         );
  AOI21_X2 U7866 ( .B1(n5851), .B2(n5850), .A(n4547), .ZN(n5852) );
  AOI21_X2 U7867 ( .B1(n4552), .B2(n5853), .A(n5852), .ZN(n5863) );
  NOR2_X4 U7868 ( .A1(n4551), .A2(n5854), .ZN(n5856) );
  MUX2_X2 U7869 ( .A(n4002), .B(n5856), .S(n5855), .Z(n5862) );
  INV_X4 U7870 ( .A(n5857), .ZN(n5860) );
  AOI221_X2 U7871 ( .B1(n5860), .B2(n8784), .C1(n4267), .C2(n5859), .A(n5858), 
        .ZN(n5861) );
  NAND3_X2 U7872 ( .A1(n5863), .A2(n5862), .A3(n5861), .ZN(out[17]) );
  NAND2_X2 U7873 ( .A1(n5864), .A2(n4401), .ZN(n5866) );
  OAI21_X4 U7874 ( .B1(n5868), .B2(n5867), .A(n5866), .ZN(n5869) );
  INV_X4 U7875 ( .A(n6072), .ZN(n5870) );
  NOR2_X4 U7876 ( .A1(n5875), .A2(n5874), .ZN(n6053) );
  NAND2_X2 U7877 ( .A1(a[15]), .A2(net246916), .ZN(n6174) );
  XOR2_X2 U7878 ( .A(n6053), .B(n6174), .Z(n5876) );
  NAND2_X2 U7879 ( .A1(a[16]), .A2(net246902), .ZN(n6052) );
  XNOR2_X2 U7880 ( .A(n5876), .B(n6052), .ZN(n6061) );
  INV_X4 U7881 ( .A(n6061), .ZN(n5883) );
  NAND2_X2 U7882 ( .A1(a[17]), .A2(n4567), .ZN(n6064) );
  INV_X4 U7883 ( .A(n6064), .ZN(n5882) );
  INV_X4 U7884 ( .A(n5877), .ZN(n5881) );
  INV_X4 U7885 ( .A(n5878), .ZN(n5880) );
  OAI21_X4 U7886 ( .B1(n5881), .B2(n5880), .A(n5879), .ZN(n6062) );
  FA_X1 U7887 ( .A(n5883), .B(n5882), .CI(n4381), .S(n6073) );
  XNOR2_X2 U7888 ( .A(n5884), .B(n6073), .ZN(n6076) );
  INV_X4 U7889 ( .A(n5885), .ZN(n5888) );
  NAND2_X2 U7890 ( .A1(n5887), .A2(n5886), .ZN(n5889) );
  NAND2_X2 U7891 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  OAI21_X4 U7892 ( .B1(n5892), .B2(n5891), .A(n5890), .ZN(n5895) );
  INV_X4 U7893 ( .A(n5895), .ZN(n5894) );
  NAND2_X2 U7894 ( .A1(a[19]), .A2(b[27]), .ZN(n5893) );
  NAND2_X2 U7895 ( .A1(a[19]), .A2(n5895), .ZN(n6194) );
  NAND2_X2 U7896 ( .A1(n6075), .A2(n6194), .ZN(n5896) );
  XNOR2_X2 U7897 ( .A(n6076), .B(n5896), .ZN(n6082) );
  INV_X4 U7898 ( .A(n6082), .ZN(n5907) );
  NAND2_X2 U7899 ( .A1(a[20]), .A2(b[26]), .ZN(n5903) );
  INV_X4 U7900 ( .A(n5903), .ZN(n5905) );
  XNOR2_X2 U7901 ( .A(n5907), .B(n5906), .ZN(n6051) );
  INV_X4 U7902 ( .A(n5911), .ZN(n6048) );
  NAND2_X2 U7903 ( .A1(n5910), .A2(n5909), .ZN(n5912) );
  INV_X4 U7904 ( .A(n5912), .ZN(n6047) );
  OAI21_X4 U7905 ( .B1(n6048), .B2(n6047), .A(a[21]), .ZN(n6049) );
  NAND2_X2 U7906 ( .A1(a[21]), .A2(b[25]), .ZN(n6045) );
  AOI21_X4 U7907 ( .B1(n5917), .B2(n5921), .A(n5916), .ZN(n5924) );
  NAND2_X2 U7908 ( .A1(a[22]), .A2(b[24]), .ZN(n5926) );
  INV_X4 U7909 ( .A(n5926), .ZN(n6088) );
  XNOR2_X2 U7910 ( .A(n5927), .B(n5928), .ZN(n5930) );
  NAND2_X2 U7911 ( .A1(net244528), .A2(net244529), .ZN(n5929) );
  XNOR2_X2 U7912 ( .A(n4010), .B(n5929), .ZN(n6031) );
  NAND2_X2 U7913 ( .A1(b[22]), .A2(a[24]), .ZN(net244537) );
  FA_X1 U7914 ( .A(n6031), .B(net244537), .CI(n5931), .S(n6023) );
  NAND2_X2 U7915 ( .A1(net246836), .A2(net246760), .ZN(n5935) );
  OAI21_X4 U7916 ( .B1(net244681), .B2(net244682), .A(net244683), .ZN(n5932)
         );
  OAI21_X4 U7917 ( .B1(n5933), .B2(net244679), .A(n5932), .ZN(n6024) );
  INV_X4 U7918 ( .A(n6024), .ZN(n5934) );
  INV_X4 U7919 ( .A(n5935), .ZN(n6025) );
  XNOR2_X2 U7920 ( .A(n6023), .B(n5936), .ZN(net244568) );
  INV_X4 U7921 ( .A(n5938), .ZN(n5941) );
  NAND2_X2 U7922 ( .A1(n5941), .A2(n5083), .ZN(n5942) );
  OAI21_X4 U7923 ( .B1(net244655), .B2(n5943), .A(n5942), .ZN(n6092) );
  XNOR2_X2 U7924 ( .A(n6093), .B(n5944), .ZN(n6098) );
  NAND2_X2 U7925 ( .A1(a[28]), .A2(b[18]), .ZN(n6096) );
  XNOR2_X2 U7926 ( .A(n5949), .B(n6096), .ZN(n5950) );
  XNOR2_X2 U7927 ( .A(n5950), .B(n6098), .ZN(n6021) );
  INV_X4 U7928 ( .A(n5954), .ZN(n5952) );
  NAND2_X2 U7929 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  INV_X4 U7930 ( .A(n5953), .ZN(n5961) );
  NAND2_X2 U7931 ( .A1(b[17]), .A2(net246788), .ZN(n5959) );
  OAI21_X4 U7932 ( .B1(n5961), .B2(n5957), .A(n5956), .ZN(n6020) );
  INV_X4 U7933 ( .A(n6020), .ZN(n5963) );
  INV_X4 U7934 ( .A(n5959), .ZN(n5960) );
  NOR3_X4 U7935 ( .A1(n5962), .A2(n5961), .A3(n5960), .ZN(n6022) );
  NOR2_X4 U7936 ( .A1(n5963), .A2(n6022), .ZN(n5964) );
  XNOR2_X2 U7937 ( .A(n5965), .B(n5964), .ZN(n6018) );
  INV_X4 U7938 ( .A(n5966), .ZN(n5967) );
  NOR3_X4 U7939 ( .A1(n5967), .A2(net247632), .A3(net244627), .ZN(n6015) );
  NAND2_X2 U7940 ( .A1(b[16]), .A2(a[30]), .ZN(n6014) );
  XNOR2_X2 U7941 ( .A(n6015), .B(n6014), .ZN(n5968) );
  XNOR2_X2 U7942 ( .A(n6018), .B(n5968), .ZN(n6107) );
  NAND2_X2 U7943 ( .A1(net240782), .A2(a[15]), .ZN(n5969) );
  NAND2_X2 U7944 ( .A1(b[15]), .A2(n5970), .ZN(n6013) );
  INV_X4 U7945 ( .A(b[15]), .ZN(net244442) );
  NAND2_X2 U7946 ( .A1(net240913), .A2(net244442), .ZN(n5971) );
  NAND2_X2 U7947 ( .A1(n5971), .A2(n4550), .ZN(n5972) );
  INV_X4 U7948 ( .A(n5973), .ZN(n5974) );
  NAND2_X2 U7949 ( .A1(n8784), .A2(n5974), .ZN(n6011) );
  NAND2_X2 U7950 ( .A1(n5976), .A2(n4579), .ZN(n5979) );
  INV_X4 U7951 ( .A(n5975), .ZN(n5978) );
  INV_X4 U7952 ( .A(n5976), .ZN(n5977) );
  AOI22_X2 U7953 ( .A1(n5979), .A2(n5978), .B1(n5977), .B2(a[16]), .ZN(n6117)
         );
  XNOR2_X2 U7954 ( .A(net246926), .B(b[15]), .ZN(n6116) );
  XNOR2_X2 U7955 ( .A(a[15]), .B(n6116), .ZN(n5980) );
  XNOR2_X2 U7956 ( .A(n6117), .B(n5980), .ZN(n6009) );
  INV_X4 U7957 ( .A(n5981), .ZN(n5984) );
  INV_X4 U7958 ( .A(n5982), .ZN(n5983) );
  OAI22_X2 U7959 ( .A1(n5984), .A2(n4539), .B1(n5983), .B2(n4531), .ZN(n6005)
         );
  AOI22_X2 U7960 ( .A1(n6564), .A2(n5985), .B1(n4557), .B2(n6280), .ZN(n5992)
         );
  INV_X4 U7961 ( .A(n8115), .ZN(n5990) );
  INV_X4 U7962 ( .A(n5986), .ZN(n5988) );
  NOR2_X4 U7963 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  OAI21_X4 U7964 ( .B1(net246956), .B2(n4580), .A(n5989), .ZN(n6920) );
  AOI22_X2 U7965 ( .A1(n5990), .A2(n6563), .B1(n6920), .B2(n4564), .ZN(n5991)
         );
  NAND2_X2 U7966 ( .A1(n5992), .A2(n5991), .ZN(n6134) );
  INV_X4 U7967 ( .A(n6134), .ZN(n5993) );
  NAND2_X2 U7968 ( .A1(n4554), .A2(n6273), .ZN(n6001) );
  NAND2_X2 U7969 ( .A1(n5994), .A2(n4565), .ZN(n6000) );
  NAND2_X2 U7970 ( .A1(net246962), .A2(a[8]), .ZN(n7038) );
  NAND2_X2 U7971 ( .A1(n4542), .A2(a[0]), .ZN(n5996) );
  NAND2_X2 U7972 ( .A1(n4562), .A2(n6913), .ZN(n5999) );
  NAND2_X2 U7973 ( .A1(n4558), .A2(n6560), .ZN(n5998) );
  NAND4_X2 U7974 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n6133)
         );
  INV_X4 U7975 ( .A(n6133), .ZN(n6002) );
  NOR3_X4 U7976 ( .A1(n6005), .A2(n6004), .A3(n6003), .ZN(n6007) );
  NAND2_X2 U7977 ( .A1(n4267), .A2(a[15]), .ZN(n6006) );
  AOI21_X2 U7978 ( .B1(n4552), .B2(n6009), .A(n6008), .ZN(n6010) );
  NAND4_X2 U7979 ( .A1(n6013), .A2(n6012), .A3(n6011), .A4(n6010), .ZN(out[15]) );
  INV_X4 U7980 ( .A(n6014), .ZN(n6016) );
  OAI21_X4 U7981 ( .B1(n6018), .B2(n6019), .A(n6017), .ZN(n6152) );
  INV_X4 U7982 ( .A(n6152), .ZN(n6155) );
  NAND2_X2 U7983 ( .A1(b[16]), .A2(net246786), .ZN(n6154) );
  INV_X4 U7984 ( .A(n6154), .ZN(n6153) );
  OAI22_X2 U7985 ( .A1(n6155), .A2(n6154), .B1(n6153), .B2(n6152), .ZN(n6106)
         );
  NAND2_X2 U7986 ( .A1(b[17]), .A2(a[28]), .ZN(n6243) );
  OAI21_X4 U7987 ( .B1(n6022), .B2(n6021), .A(n6020), .ZN(n6244) );
  XNOR2_X2 U7988 ( .A(n6243), .B(n6244), .ZN(n6104) );
  OAI21_X4 U7989 ( .B1(n6027), .B2(n6028), .A(n6026), .ZN(net244284) );
  INV_X4 U7990 ( .A(net244537), .ZN(net244545) );
  NAND2_X2 U7991 ( .A1(a[23]), .A2(b[22]), .ZN(n6033) );
  INV_X4 U7992 ( .A(n6030), .ZN(n6162) );
  INV_X4 U7993 ( .A(n6033), .ZN(n6160) );
  OAI21_X4 U7994 ( .B1(n6161), .B2(n6036), .A(n6035), .ZN(net244288) );
  INV_X4 U7995 ( .A(n6037), .ZN(n6041) );
  INV_X4 U7996 ( .A(net244529), .ZN(net244522) );
  INV_X4 U7997 ( .A(net244528), .ZN(net244523) );
  NOR3_X4 U7998 ( .A1(net244523), .A2(net244522), .A3(n6041), .ZN(n6044) );
  XNOR2_X2 U7999 ( .A(n6040), .B(n6086), .ZN(n6043) );
  OAI21_X4 U8000 ( .B1(n6044), .B2(n6043), .A(n6042), .ZN(net244369) );
  NAND2_X2 U8001 ( .A1(b[23]), .A2(a[22]), .ZN(net244371) );
  INV_X4 U8002 ( .A(n6045), .ZN(n6046) );
  NOR3_X4 U8003 ( .A1(n6048), .A2(n6047), .A3(n6046), .ZN(n6050) );
  OAI21_X4 U8004 ( .B1(n4406), .B2(n6050), .A(n6049), .ZN(n6209) );
  NAND2_X2 U8005 ( .A1(a[20]), .A2(b[25]), .ZN(n6212) );
  XNOR2_X2 U8006 ( .A(n6209), .B(n6212), .ZN(n6085) );
  NAND2_X2 U8007 ( .A1(a[14]), .A2(net249231), .ZN(n6171) );
  NAND2_X2 U8008 ( .A1(n6053), .A2(n6052), .ZN(n6055) );
  OAI21_X4 U8009 ( .B1(n6053), .B2(n6052), .A(n6174), .ZN(n6054) );
  NAND2_X2 U8010 ( .A1(n6055), .A2(n6054), .ZN(n6057) );
  INV_X4 U8011 ( .A(n6057), .ZN(n6172) );
  NAND2_X2 U8012 ( .A1(a[15]), .A2(net248516), .ZN(n6058) );
  INV_X4 U8013 ( .A(n6058), .ZN(n6056) );
  NAND2_X2 U8014 ( .A1(n6172), .A2(n6056), .ZN(n6175) );
  NAND2_X2 U8015 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  NAND2_X2 U8016 ( .A1(n6175), .A2(n6059), .ZN(n6060) );
  XNOR2_X2 U8017 ( .A(n6171), .B(n6060), .ZN(n6180) );
  INV_X4 U8018 ( .A(n6180), .ZN(n6071) );
  NAND2_X2 U8019 ( .A1(a[16]), .A2(n4567), .ZN(n6068) );
  INV_X4 U8020 ( .A(n6068), .ZN(n6066) );
  NAND2_X2 U8021 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  OAI21_X4 U8022 ( .B1(n6065), .B2(n6064), .A(n6063), .ZN(n6067) );
  NAND2_X2 U8023 ( .A1(n6066), .A2(n6067), .ZN(n6179) );
  INV_X4 U8024 ( .A(n6067), .ZN(n6069) );
  XNOR2_X2 U8025 ( .A(n6071), .B(n6070), .ZN(n6185) );
  NAND2_X2 U8026 ( .A1(a[17]), .A2(net246880), .ZN(n6187) );
  XOR2_X2 U8027 ( .A(n6185), .B(n6187), .Z(n6074) );
  OAI21_X4 U8028 ( .B1(n4439), .B2(n6073), .A(n6072), .ZN(n6184) );
  XNOR2_X2 U8029 ( .A(n6074), .B(n6184), .ZN(n6196) );
  NAND2_X2 U8030 ( .A1(n6194), .A2(n6195), .ZN(n6077) );
  XNOR2_X2 U8031 ( .A(n6196), .B(n6077), .ZN(n6079) );
  NAND2_X2 U8032 ( .A1(a[18]), .A2(b[27]), .ZN(n6199) );
  INV_X4 U8033 ( .A(n6080), .ZN(n6083) );
  OAI21_X4 U8034 ( .B1(n6083), .B2(n6082), .A(n6081), .ZN(n6165) );
  XNOR2_X2 U8035 ( .A(n4458), .B(n6165), .ZN(n6084) );
  XNOR2_X2 U8036 ( .A(n6084), .B(n3935), .ZN(n6208) );
  XNOR2_X2 U8037 ( .A(n6085), .B(n4446), .ZN(n6220) );
  NAND2_X2 U8038 ( .A1(a[21]), .A2(b[24]), .ZN(n6221) );
  XNOR2_X2 U8039 ( .A(n6219), .B(n6221), .ZN(n6089) );
  XNOR2_X2 U8040 ( .A(n6224), .B(n6089), .ZN(net244368) );
  AOI21_X4 U8041 ( .B1(n3965), .B2(n6093), .A(n6091), .ZN(n6095) );
  NAND2_X2 U8042 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  XNOR2_X2 U8043 ( .A(net244457), .B(net247881), .ZN(net244258) );
  NAND2_X2 U8044 ( .A1(b[18]), .A2(net246772), .ZN(net244260) );
  INV_X4 U8045 ( .A(n6096), .ZN(n6100) );
  OAI21_X4 U8046 ( .B1(n6099), .B2(n6100), .A(n6098), .ZN(n6241) );
  XNOR2_X2 U8047 ( .A(n6102), .B(net244258), .ZN(n6311) );
  INV_X4 U8048 ( .A(n6311), .ZN(n6103) );
  XNOR2_X2 U8049 ( .A(n6104), .B(n6103), .ZN(n6156) );
  XNOR2_X2 U8050 ( .A(n6106), .B(n6105), .ZN(n6150) );
  INV_X4 U8051 ( .A(n6107), .ZN(n6108) );
  NOR3_X4 U8052 ( .A1(n6108), .A2(net246812), .A3(net244442), .ZN(n6147) );
  NAND2_X2 U8053 ( .A1(b[15]), .A2(a[30]), .ZN(n6146) );
  XNOR2_X2 U8054 ( .A(n6147), .B(n6146), .ZN(n6109) );
  XNOR2_X2 U8055 ( .A(n6150), .B(n6109), .ZN(n6255) );
  NAND2_X2 U8056 ( .A1(net240782), .A2(a[14]), .ZN(n6110) );
  NAND2_X2 U8057 ( .A1(b[14]), .A2(n6111), .ZN(n6145) );
  NAND2_X2 U8058 ( .A1(net240913), .A2(net244239), .ZN(n6112) );
  NAND2_X2 U8059 ( .A1(n6112), .A2(n4550), .ZN(n6113) );
  INV_X4 U8060 ( .A(n6114), .ZN(n6115) );
  NAND2_X2 U8061 ( .A1(n8784), .A2(n6115), .ZN(n6143) );
  XNOR2_X2 U8062 ( .A(net246926), .B(b[14]), .ZN(n6264) );
  XNOR2_X2 U8063 ( .A(a[14]), .B(n6264), .ZN(n6121) );
  INV_X4 U8064 ( .A(n6116), .ZN(n6119) );
  NAND2_X2 U8065 ( .A1(n6117), .A2(n4580), .ZN(n6118) );
  OAI21_X4 U8066 ( .B1(n6120), .B2(n6119), .A(n6118), .ZN(n6265) );
  XNOR2_X2 U8067 ( .A(n6121), .B(n6265), .ZN(n6141) );
  NOR2_X4 U8068 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  OAI21_X4 U8069 ( .B1(net246956), .B2(n4581), .A(n6126), .ZN(n7039) );
  AOI22_X2 U8070 ( .A1(n7039), .A2(n4564), .B1(n4555), .B2(n6699), .ZN(n6127)
         );
  NAND2_X2 U8071 ( .A1(n6128), .A2(n6127), .ZN(n6270) );
  INV_X4 U8072 ( .A(n6270), .ZN(n6136) );
  INV_X4 U8073 ( .A(n6697), .ZN(n6131) );
  AOI22_X2 U8074 ( .A1(n6129), .A2(n4565), .B1(n4555), .B2(n6404), .ZN(n6130)
         );
  OAI221_X2 U8075 ( .B1(n6131), .B2(n8832), .C1(n853), .C2(n4533), .A(n6130), 
        .ZN(n6132) );
  INV_X4 U8076 ( .A(n6132), .ZN(n6272) );
  AOI22_X2 U8077 ( .A1(n8841), .A2(n6134), .B1(n8842), .B2(n6133), .ZN(n6135)
         );
  OAI221_X2 U8078 ( .B1(n6136), .B2(n4537), .C1(n6272), .C2(n4535), .A(n6135), 
        .ZN(n6137) );
  INV_X4 U8079 ( .A(n6137), .ZN(n6139) );
  NAND2_X2 U8080 ( .A1(net247002), .A2(a[14]), .ZN(n6138) );
  AOI21_X2 U8081 ( .B1(n4552), .B2(n6141), .A(n6140), .ZN(n6142) );
  NAND4_X2 U8082 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(out[14]) );
  INV_X4 U8083 ( .A(n6146), .ZN(n6148) );
  OAI21_X4 U8084 ( .B1(n6150), .B2(n6151), .A(n6149), .ZN(n6383) );
  INV_X4 U8085 ( .A(n6383), .ZN(n6382) );
  NAND2_X2 U8086 ( .A1(b[15]), .A2(net246788), .ZN(n6381) );
  INV_X4 U8087 ( .A(n6381), .ZN(n6384) );
  NAND2_X2 U8088 ( .A1(a[28]), .A2(b[16]), .ZN(n6307) );
  INV_X4 U8089 ( .A(n6307), .ZN(n6159) );
  NAND2_X2 U8090 ( .A1(n6155), .A2(n6154), .ZN(n6157) );
  NAND2_X2 U8091 ( .A1(n6157), .A2(n6156), .ZN(n6305) );
  XNOR2_X2 U8092 ( .A(n6159), .B(n6158), .ZN(n6253) );
  XOR2_X2 U8093 ( .A(net244136), .B(n6322), .Z(n6235) );
  INV_X4 U8094 ( .A(net244371), .ZN(net244370) );
  INV_X4 U8095 ( .A(n6326), .ZN(n6164) );
  NAND2_X2 U8096 ( .A1(a[21]), .A2(b[23]), .ZN(n6330) );
  NAND3_X2 U8097 ( .A1(n6329), .A2(n6328), .A3(n6330), .ZN(n6163) );
  OAI21_X4 U8098 ( .B1(n6164), .B2(n4572), .A(n6163), .ZN(n6234) );
  OAI21_X4 U8099 ( .B1(n4457), .B2(n6166), .A(n3935), .ZN(n6168) );
  NAND2_X2 U8100 ( .A1(n6166), .A2(n4458), .ZN(n6167) );
  AOI21_X4 U8101 ( .B1(a[18]), .B2(b[26]), .A(n6169), .ZN(n6336) );
  NAND2_X2 U8102 ( .A1(a[18]), .A2(n6169), .ZN(n6334) );
  INV_X4 U8103 ( .A(n6334), .ZN(n6170) );
  INV_X4 U8104 ( .A(n6171), .ZN(n6173) );
  NAND2_X2 U8105 ( .A1(n6173), .A2(n6172), .ZN(n6176) );
  NAND2_X2 U8106 ( .A1(a[14]), .A2(net248517), .ZN(n6341) );
  NAND3_X2 U8107 ( .A1(n6176), .A2(n6175), .A3(n3962), .ZN(n6342) );
  NAND2_X2 U8108 ( .A1(a[13]), .A2(net246916), .ZN(n6446) );
  XNOR2_X2 U8109 ( .A(n6341), .B(n6446), .ZN(n6177) );
  XNOR2_X2 U8110 ( .A(n6342), .B(n6177), .ZN(n6347) );
  INV_X4 U8111 ( .A(n6347), .ZN(n6183) );
  NAND2_X2 U8112 ( .A1(a[15]), .A2(n4567), .ZN(n6350) );
  INV_X4 U8113 ( .A(n6350), .ZN(n6182) );
  INV_X4 U8114 ( .A(n6178), .ZN(n6181) );
  OAI21_X4 U8115 ( .B1(n6181), .B2(n6180), .A(n6179), .ZN(n6348) );
  FA_X1 U8116 ( .A(n6183), .B(n6182), .CI(n6348), .S(n6360) );
  NAND2_X2 U8117 ( .A1(a[16]), .A2(net246880), .ZN(n6191) );
  INV_X4 U8118 ( .A(n6191), .ZN(n6189) );
  NAND2_X2 U8119 ( .A1(n6189), .A2(n6190), .ZN(n6359) );
  INV_X4 U8120 ( .A(n6190), .ZN(n6192) );
  XNOR2_X2 U8121 ( .A(n6360), .B(n6193), .ZN(n6339) );
  NAND2_X2 U8122 ( .A1(a[17]), .A2(b[27]), .ZN(n6203) );
  INV_X4 U8123 ( .A(n6203), .ZN(n6201) );
  NAND2_X2 U8124 ( .A1(n6195), .A2(n6194), .ZN(n6197) );
  NAND2_X2 U8125 ( .A1(n6197), .A2(n6196), .ZN(n6198) );
  OAI21_X4 U8126 ( .B1(n6200), .B2(n6199), .A(n6198), .ZN(n6202) );
  NAND2_X2 U8127 ( .A1(n6201), .A2(n6202), .ZN(n6338) );
  INV_X4 U8128 ( .A(n6202), .ZN(n6204) );
  NAND2_X2 U8129 ( .A1(n6204), .A2(n6203), .ZN(n6337) );
  NAND2_X2 U8130 ( .A1(n6338), .A2(n6337), .ZN(n6205) );
  XNOR2_X2 U8131 ( .A(n6339), .B(n6205), .ZN(n6335) );
  INV_X4 U8132 ( .A(n6335), .ZN(n6206) );
  XNOR2_X2 U8133 ( .A(n6207), .B(n6206), .ZN(n6367) );
  NAND2_X2 U8134 ( .A1(a[19]), .A2(b[25]), .ZN(n6216) );
  INV_X4 U8135 ( .A(n6216), .ZN(n6214) );
  INV_X4 U8136 ( .A(n6208), .ZN(n6210) );
  OAI21_X4 U8137 ( .B1(n6213), .B2(n6212), .A(n6211), .ZN(n6215) );
  NAND2_X2 U8138 ( .A1(n6214), .A2(n6215), .ZN(n6366) );
  INV_X4 U8139 ( .A(n6215), .ZN(n6217) );
  NAND2_X2 U8140 ( .A1(n6366), .A2(n6365), .ZN(n6218) );
  XNOR2_X2 U8141 ( .A(n6367), .B(n6218), .ZN(n6371) );
  NAND2_X2 U8142 ( .A1(n6220), .A2(n6219), .ZN(n6231) );
  INV_X4 U8143 ( .A(n6231), .ZN(n6229) );
  INV_X4 U8144 ( .A(n6221), .ZN(n6226) );
  INV_X4 U8145 ( .A(n6230), .ZN(n6228) );
  NAND2_X2 U8146 ( .A1(a[20]), .A2(b[24]), .ZN(n6232) );
  INV_X4 U8147 ( .A(n6232), .ZN(n6227) );
  OAI21_X4 U8148 ( .B1(n6229), .B2(n6228), .A(n6227), .ZN(n6370) );
  NAND3_X4 U8149 ( .A1(n6230), .A2(n6231), .A3(n6232), .ZN(n6495) );
  NAND2_X2 U8150 ( .A1(n6370), .A2(n6495), .ZN(n6233) );
  XNOR2_X2 U8151 ( .A(n6233), .B(n6371), .ZN(n6327) );
  XNOR2_X2 U8152 ( .A(n6234), .B(n4391), .ZN(n6321) );
  XNOR2_X2 U8153 ( .A(n6235), .B(n6321), .ZN(n6320) );
  INV_X4 U8154 ( .A(net244283), .ZN(net244287) );
  NAND2_X2 U8155 ( .A1(net244283), .A2(net244284), .ZN(net244145) );
  NAND2_X2 U8156 ( .A1(net246836), .A2(a[23]), .ZN(n6316) );
  XNOR2_X2 U8157 ( .A(n6239), .B(n6238), .ZN(net244075) );
  NAND2_X2 U8158 ( .A1(b[20]), .A2(a[24]), .ZN(net244078) );
  XNOR2_X2 U8159 ( .A(net244256), .B(net244257), .ZN(n6246) );
  NAND2_X2 U8160 ( .A1(n6242), .A2(n6243), .ZN(n6310) );
  NAND2_X2 U8161 ( .A1(b[17]), .A2(net246772), .ZN(n6248) );
  INV_X4 U8162 ( .A(n6243), .ZN(n6245) );
  INV_X4 U8163 ( .A(n6248), .ZN(n6314) );
  NAND3_X2 U8164 ( .A1(n6246), .A2(n6310), .A3(n6314), .ZN(n6247) );
  INV_X4 U8165 ( .A(n6247), .ZN(n6250) );
  NOR3_X4 U8166 ( .A1(n6251), .A2(n6250), .A3(n6249), .ZN(n6252) );
  XNOR2_X2 U8167 ( .A(net244244), .B(n6252), .ZN(net244177) );
  INV_X4 U8168 ( .A(net244177), .ZN(net244243) );
  XNOR2_X2 U8169 ( .A(n4422), .B(net244243), .ZN(n6428) );
  XNOR2_X2 U8170 ( .A(n4464), .B(n6254), .ZN(n6302) );
  INV_X4 U8171 ( .A(n6255), .ZN(n6256) );
  NOR3_X4 U8172 ( .A1(n6256), .A2(net247632), .A3(net244239), .ZN(n6299) );
  NAND2_X2 U8173 ( .A1(b[14]), .A2(a[30]), .ZN(n6298) );
  XNOR2_X2 U8174 ( .A(n6299), .B(n6298), .ZN(n6257) );
  NAND2_X2 U8175 ( .A1(net240782), .A2(a[13]), .ZN(n6258) );
  NAND2_X2 U8176 ( .A1(b[13]), .A2(n6259), .ZN(n6297) );
  NAND2_X2 U8177 ( .A1(net240913), .A2(n6389), .ZN(n6260) );
  NAND2_X2 U8178 ( .A1(n6260), .A2(n4550), .ZN(n6261) );
  INV_X4 U8179 ( .A(n6262), .ZN(n6263) );
  NAND2_X2 U8180 ( .A1(n8784), .A2(n6263), .ZN(n6295) );
  NAND2_X2 U8181 ( .A1(n6265), .A2(n4581), .ZN(n6268) );
  INV_X4 U8182 ( .A(n6264), .ZN(n6267) );
  INV_X4 U8183 ( .A(n6265), .ZN(n6266) );
  AOI22_X2 U8184 ( .A1(n6268), .A2(n6267), .B1(n6266), .B2(a[14]), .ZN(n6399)
         );
  XNOR2_X2 U8185 ( .A(net246924), .B(b[13]), .ZN(n6397) );
  XNOR2_X2 U8186 ( .A(a[13]), .B(n6397), .ZN(n6269) );
  XNOR2_X2 U8187 ( .A(n6399), .B(n6269), .ZN(n6293) );
  NAND2_X2 U8188 ( .A1(n8841), .A2(n6270), .ZN(n6271) );
  INV_X4 U8189 ( .A(n6913), .ZN(n6276) );
  NAND2_X2 U8190 ( .A1(n7044), .A2(n3982), .ZN(n7256) );
  INV_X4 U8191 ( .A(n7256), .ZN(n6275) );
  AOI22_X2 U8192 ( .A1(n6273), .A2(n4565), .B1(n4554), .B2(n6560), .ZN(n6274)
         );
  OAI221_X2 U8193 ( .B1(n6276), .B2(n8832), .C1(n6275), .C2(n4533), .A(n6274), 
        .ZN(n6277) );
  INV_X4 U8194 ( .A(n6277), .ZN(n6418) );
  INV_X4 U8195 ( .A(n6563), .ZN(n6278) );
  NAND2_X2 U8196 ( .A1(net247082), .A2(net246790), .ZN(n6281) );
  AOI22_X2 U8197 ( .A1(n4555), .A2(n6920), .B1(n7247), .B2(n4564), .ZN(n6284)
         );
  NAND2_X2 U8198 ( .A1(n6285), .A2(n6284), .ZN(n6416) );
  INV_X4 U8199 ( .A(n6416), .ZN(n6286) );
  NOR3_X4 U8200 ( .A1(n6289), .A2(n6288), .A3(n6287), .ZN(n6291) );
  NAND2_X2 U8201 ( .A1(net247002), .A2(a[13]), .ZN(n6290) );
  AOI21_X2 U8202 ( .B1(n4552), .B2(n6293), .A(n6292), .ZN(n6294) );
  NAND4_X2 U8203 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(out[13]) );
  INV_X4 U8204 ( .A(n6298), .ZN(n6300) );
  OAI21_X4 U8205 ( .B1(n6303), .B2(n6302), .A(n6301), .ZN(n6535) );
  NAND2_X2 U8206 ( .A1(b[14]), .A2(net246788), .ZN(n6531) );
  INV_X4 U8207 ( .A(n6531), .ZN(n6536) );
  OAI22_X2 U8208 ( .A1(n6532), .A2(n6531), .B1(n6536), .B2(n6535), .ZN(n6387)
         );
  NAND2_X2 U8209 ( .A1(n6305), .A2(n6304), .ZN(n6308) );
  INV_X4 U8210 ( .A(n6308), .ZN(n6306) );
  NAND2_X2 U8211 ( .A1(n6306), .A2(n6307), .ZN(net244178) );
  NAND2_X2 U8212 ( .A1(net244177), .A2(net244178), .ZN(n6309) );
  NAND2_X2 U8213 ( .A1(n6159), .A2(n6308), .ZN(net244181) );
  NAND2_X2 U8214 ( .A1(b[16]), .A2(net246772), .ZN(net244180) );
  OAI21_X4 U8215 ( .B1(n6315), .B2(n3906), .A(n6314), .ZN(n6529) );
  XNOR2_X2 U8216 ( .A(net243763), .B(net243760), .ZN(net244064) );
  NAND2_X2 U8217 ( .A1(net246760), .A2(b[18]), .ZN(net244156) );
  INV_X4 U8218 ( .A(n6316), .ZN(n6317) );
  NAND2_X2 U8219 ( .A1(net246836), .A2(a[22]), .ZN(n6441) );
  XOR2_X2 U8220 ( .A(n6438), .B(n6441), .Z(n6376) );
  INV_X4 U8221 ( .A(n6321), .ZN(n6323) );
  INV_X4 U8222 ( .A(n6322), .ZN(n6324) );
  OAI21_X4 U8223 ( .B1(n6323), .B2(n6324), .A(net244136), .ZN(n6520) );
  XNOR2_X2 U8224 ( .A(n3939), .B(n6325), .ZN(n6375) );
  NAND2_X2 U8225 ( .A1(a[21]), .A2(n6326), .ZN(n6508) );
  INV_X4 U8226 ( .A(n6327), .ZN(n6332) );
  NAND2_X2 U8227 ( .A1(n6507), .A2(n6508), .ZN(n6333) );
  NAND2_X2 U8228 ( .A1(a[20]), .A2(b[23]), .ZN(n6512) );
  XNOR2_X2 U8229 ( .A(n6333), .B(n6512), .ZN(n6373) );
  NAND2_X2 U8230 ( .A1(a[19]), .A2(b[24]), .ZN(n6500) );
  OAI21_X4 U8231 ( .B1(n6336), .B2(n6335), .A(n6334), .ZN(n6477) );
  NAND2_X2 U8232 ( .A1(a[17]), .A2(b[26]), .ZN(n6475) );
  INV_X4 U8233 ( .A(n6337), .ZN(n6340) );
  NAND2_X2 U8234 ( .A1(a[15]), .A2(net246880), .ZN(n6458) );
  NAND2_X2 U8235 ( .A1(a[12]), .A2(net249231), .ZN(n6444) );
  INV_X4 U8236 ( .A(n6341), .ZN(n6343) );
  NAND2_X2 U8237 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  OAI21_X4 U8238 ( .B1(n6345), .B2(n6446), .A(n6344), .ZN(n6443) );
  XOR2_X2 U8239 ( .A(n6444), .B(n6443), .Z(n6346) );
  NAND2_X2 U8240 ( .A1(a[13]), .A2(net246902), .ZN(n6445) );
  XNOR2_X2 U8241 ( .A(n6346), .B(n6445), .ZN(n6451) );
  INV_X4 U8242 ( .A(n6451), .ZN(n6357) );
  NAND2_X2 U8243 ( .A1(a[14]), .A2(n4567), .ZN(n6354) );
  INV_X4 U8244 ( .A(n6354), .ZN(n6352) );
  NAND2_X2 U8245 ( .A1(n6348), .A2(n6347), .ZN(n6349) );
  OAI21_X4 U8246 ( .B1(n6351), .B2(n6350), .A(n6349), .ZN(n6353) );
  NAND2_X2 U8247 ( .A1(n6352), .A2(n6353), .ZN(n6450) );
  INV_X4 U8248 ( .A(n6353), .ZN(n6355) );
  NAND2_X2 U8249 ( .A1(n6355), .A2(n6354), .ZN(n6449) );
  NAND2_X2 U8250 ( .A1(n6450), .A2(n6449), .ZN(n6356) );
  XNOR2_X2 U8251 ( .A(n6357), .B(n6356), .ZN(n6456) );
  INV_X4 U8252 ( .A(n6358), .ZN(n6361) );
  OAI21_X4 U8253 ( .B1(n6361), .B2(n6360), .A(n6359), .ZN(n6455) );
  XNOR2_X2 U8254 ( .A(n6455), .B(n6456), .ZN(n6362) );
  XNOR2_X2 U8255 ( .A(n6362), .B(n6458), .ZN(n6465) );
  INV_X4 U8256 ( .A(n6365), .ZN(n6368) );
  OAI21_X4 U8257 ( .B1(n6368), .B2(n6367), .A(n6366), .ZN(n6485) );
  XNOR2_X2 U8258 ( .A(n6369), .B(n3969), .ZN(n6497) );
  XNOR2_X2 U8259 ( .A(n6497), .B(n6496), .ZN(n6372) );
  XNOR2_X2 U8260 ( .A(n6500), .B(n6372), .ZN(n6510) );
  XNOR2_X2 U8261 ( .A(n6373), .B(n6510), .ZN(n6374) );
  INV_X4 U8262 ( .A(n6374), .ZN(n6521) );
  XNOR2_X2 U8263 ( .A(n6375), .B(n6521), .ZN(n6439) );
  XNOR2_X2 U8264 ( .A(n6376), .B(n6439), .ZN(n6432) );
  INV_X4 U8265 ( .A(n6432), .ZN(n6380) );
  NAND2_X2 U8266 ( .A1(a[23]), .A2(b[20]), .ZN(n6378) );
  INV_X4 U8267 ( .A(n6378), .ZN(n6434) );
  OAI22_X2 U8268 ( .A1(n6378), .A2(n6377), .B1(n6434), .B2(n6433), .ZN(n6379)
         );
  XNOR2_X2 U8269 ( .A(n6379), .B(n6380), .ZN(net243991) );
  NAND2_X2 U8270 ( .A1(b[15]), .A2(a[28]), .ZN(net244008) );
  INV_X4 U8271 ( .A(n6430), .ZN(n6385) );
  XNOR2_X2 U8272 ( .A(n6386), .B(n6387), .ZN(n6542) );
  NOR3_X4 U8273 ( .A1(n4434), .A2(net246812), .A3(n6389), .ZN(n6539) );
  NAND2_X2 U8274 ( .A1(b[13]), .A2(a[30]), .ZN(n6538) );
  XNOR2_X2 U8275 ( .A(n6539), .B(n6538), .ZN(n6390) );
  XNOR2_X2 U8276 ( .A(n6542), .B(n6390), .ZN(n6545) );
  NAND2_X2 U8277 ( .A1(net240782), .A2(a[12]), .ZN(n6391) );
  NAND2_X2 U8278 ( .A1(b[12]), .A2(n6392), .ZN(n6427) );
  NAND2_X2 U8279 ( .A1(net240913), .A2(net243844), .ZN(n6393) );
  NAND2_X2 U8280 ( .A1(n6393), .A2(n4550), .ZN(n6394) );
  INV_X4 U8281 ( .A(n6395), .ZN(n6396) );
  NAND2_X2 U8282 ( .A1(n8784), .A2(n6396), .ZN(n6425) );
  XNOR2_X2 U8283 ( .A(net246924), .B(b[12]), .ZN(n6554) );
  XNOR2_X2 U8284 ( .A(a[12]), .B(n6554), .ZN(n6403) );
  INV_X4 U8285 ( .A(n6397), .ZN(n6401) );
  NAND2_X2 U8286 ( .A1(n6399), .A2(n6398), .ZN(n6400) );
  OAI21_X4 U8287 ( .B1(n6402), .B2(n6401), .A(n6400), .ZN(n6555) );
  XNOR2_X2 U8288 ( .A(n6403), .B(n6555), .ZN(n6423) );
  INV_X4 U8289 ( .A(n7415), .ZN(n6406) );
  AOI22_X2 U8290 ( .A1(n6404), .A2(n4565), .B1(n4554), .B2(n6697), .ZN(n6405)
         );
  OAI221_X2 U8291 ( .B1(n6406), .B2(n4533), .C1(n853), .C2(n8832), .A(n6405), 
        .ZN(n6407) );
  INV_X4 U8292 ( .A(n6407), .ZN(n6574) );
  NAND2_X2 U8293 ( .A1(n4554), .A2(n7039), .ZN(n6415) );
  NAND2_X2 U8294 ( .A1(n4562), .A2(n6408), .ZN(n6414) );
  NAND2_X2 U8295 ( .A1(net247082), .A2(a[28]), .ZN(n6409) );
  NAND2_X2 U8296 ( .A1(n7419), .A2(n4565), .ZN(n6413) );
  NAND2_X2 U8297 ( .A1(n4558), .A2(n6699), .ZN(n6412) );
  NAND4_X2 U8298 ( .A1(n6415), .A2(n6414), .A3(n6413), .A4(n6412), .ZN(n6572)
         );
  AOI22_X2 U8299 ( .A1(n8318), .A2(n6572), .B1(n8841), .B2(n6416), .ZN(n6417)
         );
  OAI221_X2 U8300 ( .B1(n6418), .B2(n4531), .C1(n6574), .C2(n4535), .A(n6417), 
        .ZN(n6419) );
  INV_X4 U8301 ( .A(n6419), .ZN(n6421) );
  NAND2_X2 U8302 ( .A1(net247002), .A2(a[12]), .ZN(n6420) );
  AOI21_X2 U8303 ( .B1(n4552), .B2(n6423), .A(n6422), .ZN(n6424) );
  NAND4_X2 U8304 ( .A1(n6427), .A2(n6426), .A3(n6425), .A4(n6424), .ZN(out[12]) );
  INV_X4 U8305 ( .A(n6428), .ZN(n6429) );
  NAND3_X2 U8306 ( .A1(net244005), .A2(net244006), .A3(net244008), .ZN(n6431)
         );
  NAND2_X2 U8307 ( .A1(net243999), .A2(n6431), .ZN(net243785) );
  NAND2_X2 U8308 ( .A1(b[19]), .A2(a[23]), .ZN(net243733) );
  NAND2_X2 U8309 ( .A1(a[22]), .A2(b[20]), .ZN(n6672) );
  XNOR2_X2 U8310 ( .A(n6674), .B(n6672), .ZN(n6528) );
  NAND2_X2 U8311 ( .A1(n6439), .A2(n4466), .ZN(n6440) );
  OAI21_X4 U8312 ( .B1(n6442), .B2(n6441), .A(n6440), .ZN(n6746) );
  INV_X4 U8313 ( .A(n6443), .ZN(n6447) );
  NAND2_X2 U8314 ( .A1(a[12]), .A2(net246904), .ZN(n6624) );
  OAI21_X4 U8315 ( .B1(n6447), .B2(n3936), .A(n3961), .ZN(n6625) );
  NAND2_X2 U8316 ( .A1(a[11]), .A2(net246916), .ZN(n6628) );
  XNOR2_X2 U8317 ( .A(n6624), .B(n6628), .ZN(n6448) );
  XNOR2_X2 U8318 ( .A(n6625), .B(n6448), .ZN(n6632) );
  INV_X4 U8319 ( .A(n6632), .ZN(n6454) );
  NAND2_X2 U8320 ( .A1(a[13]), .A2(b[29]), .ZN(n6635) );
  INV_X4 U8321 ( .A(n6635), .ZN(n6453) );
  INV_X4 U8322 ( .A(n6449), .ZN(n6452) );
  OAI21_X4 U8323 ( .B1(n6452), .B2(n6451), .A(n6450), .ZN(n6633) );
  FA_X1 U8324 ( .A(n6454), .B(n6453), .CI(n6633), .S(n6622) );
  NAND2_X2 U8325 ( .A1(a[14]), .A2(net246880), .ZN(n6462) );
  INV_X4 U8326 ( .A(n6462), .ZN(n6460) );
  OAI21_X4 U8327 ( .B1(n6459), .B2(n6458), .A(n6457), .ZN(n6461) );
  INV_X4 U8328 ( .A(n6461), .ZN(n6463) );
  NAND2_X2 U8329 ( .A1(n6463), .A2(n6462), .ZN(n6620) );
  NAND2_X2 U8330 ( .A1(n6621), .A2(n6620), .ZN(n6464) );
  XNOR2_X2 U8331 ( .A(n6622), .B(n6464), .ZN(n6618) );
  NAND2_X2 U8332 ( .A1(n6466), .A2(n6467), .ZN(n6472) );
  OAI21_X4 U8333 ( .B1(n6467), .B2(n6466), .A(n3968), .ZN(n6471) );
  NAND2_X2 U8334 ( .A1(a[15]), .A2(b[27]), .ZN(n6473) );
  INV_X4 U8335 ( .A(n6473), .ZN(n6468) );
  OAI21_X4 U8336 ( .B1(n6470), .B2(n6469), .A(n6468), .ZN(n6617) );
  XNOR2_X2 U8337 ( .A(n6618), .B(n6474), .ZN(n6647) );
  INV_X4 U8338 ( .A(n6482), .ZN(n6480) );
  INV_X4 U8339 ( .A(n6475), .ZN(n6476) );
  OAI21_X4 U8340 ( .B1(n4470), .B2(n6477), .A(n6476), .ZN(n6481) );
  NAND2_X2 U8341 ( .A1(a[16]), .A2(b[26]), .ZN(n6483) );
  INV_X4 U8342 ( .A(n6483), .ZN(n6478) );
  OAI21_X4 U8343 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(n6646) );
  NAND3_X4 U8344 ( .A1(n6483), .A2(n6482), .A3(n6481), .ZN(n6645) );
  NAND2_X2 U8345 ( .A1(n4454), .A2(n6645), .ZN(n6484) );
  XNOR2_X2 U8346 ( .A(n6647), .B(n6484), .ZN(n6651) );
  NAND2_X2 U8347 ( .A1(a[17]), .A2(b[25]), .ZN(n6491) );
  INV_X4 U8348 ( .A(n6491), .ZN(n6489) );
  NAND2_X2 U8349 ( .A1(n6489), .A2(n6490), .ZN(n6650) );
  XNOR2_X2 U8350 ( .A(n4372), .B(n6493), .ZN(n6614) );
  NAND2_X2 U8351 ( .A1(a[18]), .A2(b[24]), .ZN(n6504) );
  INV_X4 U8352 ( .A(n6504), .ZN(n6502) );
  INV_X4 U8353 ( .A(n6496), .ZN(n6498) );
  NAND2_X2 U8354 ( .A1(n6498), .A2(n6497), .ZN(n6499) );
  OAI21_X4 U8355 ( .B1(n6501), .B2(n6500), .A(n6499), .ZN(n6503) );
  NAND2_X2 U8356 ( .A1(n6502), .A2(n6503), .ZN(n6613) );
  INV_X4 U8357 ( .A(n6503), .ZN(n6505) );
  NAND2_X2 U8358 ( .A1(n6505), .A2(n6504), .ZN(n6612) );
  NAND2_X2 U8359 ( .A1(n6613), .A2(n6612), .ZN(n6506) );
  XNOR2_X2 U8360 ( .A(n6614), .B(n6506), .ZN(n6657) );
  NAND2_X2 U8361 ( .A1(a[19]), .A2(b[23]), .ZN(n6516) );
  INV_X4 U8362 ( .A(n6516), .ZN(n6514) );
  NAND2_X2 U8363 ( .A1(n6510), .A2(n6509), .ZN(n6511) );
  OAI21_X4 U8364 ( .B1(n6513), .B2(n6512), .A(n6511), .ZN(n6515) );
  NAND2_X2 U8365 ( .A1(n6514), .A2(n6515), .ZN(n6656) );
  INV_X4 U8366 ( .A(n6515), .ZN(n6517) );
  NAND2_X2 U8367 ( .A1(n6656), .A2(n6655), .ZN(n6518) );
  XNOR2_X2 U8368 ( .A(n6657), .B(n6518), .ZN(n6662) );
  NAND2_X2 U8369 ( .A1(a[20]), .A2(b[22]), .ZN(n6524) );
  INV_X4 U8370 ( .A(n6524), .ZN(n6525) );
  OAI21_X4 U8371 ( .B1(n6521), .B2(n6325), .A(n3939), .ZN(n6523) );
  NAND2_X2 U8372 ( .A1(n6325), .A2(n6521), .ZN(n6522) );
  XNOR2_X2 U8373 ( .A(n6662), .B(n6526), .ZN(n6666) );
  XNOR2_X2 U8374 ( .A(n6527), .B(n4418), .ZN(n6673) );
  XNOR2_X2 U8375 ( .A(n6528), .B(n6673), .ZN(net243723) );
  NAND2_X2 U8376 ( .A1(b[17]), .A2(net246760), .ZN(net243761) );
  INV_X4 U8377 ( .A(n6683), .ZN(n6681) );
  XNOR2_X2 U8378 ( .A(net243639), .B(n6681), .ZN(n6537) );
  NAND2_X2 U8379 ( .A1(n6532), .A2(n6531), .ZN(n6534) );
  XNOR2_X2 U8380 ( .A(n6537), .B(n6682), .ZN(n6884) );
  INV_X4 U8381 ( .A(n6538), .ZN(n6540) );
  NAND2_X2 U8382 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  OAI21_X4 U8383 ( .B1(n6542), .B2(n6543), .A(n6541), .ZN(n6591) );
  INV_X4 U8384 ( .A(n6591), .ZN(n6594) );
  NAND2_X2 U8385 ( .A1(b[13]), .A2(net246790), .ZN(n6593) );
  INV_X4 U8386 ( .A(n6593), .ZN(n6592) );
  XNOR2_X2 U8387 ( .A(n6596), .B(n6544), .ZN(n6589) );
  INV_X4 U8388 ( .A(n6545), .ZN(n6546) );
  NOR3_X4 U8389 ( .A1(n6546), .A2(net247632), .A3(net243844), .ZN(n6586) );
  NAND2_X2 U8390 ( .A1(b[12]), .A2(a[30]), .ZN(n6585) );
  XNOR2_X2 U8391 ( .A(n6586), .B(n6585), .ZN(n6547) );
  XNOR2_X2 U8392 ( .A(n4436), .B(n6547), .ZN(n6687) );
  NAND2_X2 U8393 ( .A1(net240782), .A2(a[11]), .ZN(n6548) );
  NAND2_X2 U8394 ( .A1(b[11]), .A2(n6549), .ZN(n6584) );
  NAND2_X2 U8395 ( .A1(net240913), .A2(net243628), .ZN(n6550) );
  NAND2_X2 U8396 ( .A1(n6550), .A2(n4550), .ZN(n6551) );
  NAND2_X2 U8397 ( .A1(n8784), .A2(n6552), .ZN(n6582) );
  NAND2_X2 U8398 ( .A1(n6555), .A2(n6553), .ZN(n6558) );
  INV_X4 U8399 ( .A(n6554), .ZN(n6557) );
  INV_X4 U8400 ( .A(n6555), .ZN(n6556) );
  AOI22_X2 U8401 ( .A1(n6558), .A2(n6557), .B1(n6556), .B2(a[12]), .ZN(n6713)
         );
  XNOR2_X2 U8402 ( .A(net246924), .B(b[11]), .ZN(n6711) );
  XNOR2_X2 U8403 ( .A(a[11]), .B(n6711), .ZN(n6559) );
  XNOR2_X2 U8404 ( .A(n6713), .B(n6559), .ZN(n6580) );
  NAND2_X2 U8405 ( .A1(n4558), .A2(n7256), .ZN(n6562) );
  AOI22_X2 U8406 ( .A1(n6560), .A2(n4565), .B1(n4554), .B2(n6913), .ZN(n6561)
         );
  OAI211_X2 U8407 ( .C1(n949), .C2(n4533), .A(n6562), .B(n6561), .ZN(n6696) );
  INV_X4 U8408 ( .A(n6696), .ZN(n6571) );
  NAND2_X2 U8409 ( .A1(n4558), .A2(n6920), .ZN(n6569) );
  NAND2_X2 U8410 ( .A1(n6564), .A2(n6563), .ZN(n6568) );
  NAND2_X2 U8411 ( .A1(n4554), .A2(n7247), .ZN(n6567) );
  NAND2_X2 U8412 ( .A1(n7658), .A2(n4565), .ZN(n6566) );
  NAND4_X2 U8413 ( .A1(n6569), .A2(n6568), .A3(n6567), .A4(n6566), .ZN(n6693)
         );
  NAND2_X2 U8414 ( .A1(n8318), .A2(n6693), .ZN(n6570) );
  NAND2_X2 U8415 ( .A1(n8841), .A2(n6572), .ZN(n6573) );
  NOR2_X4 U8416 ( .A1(n6576), .A2(n6575), .ZN(n6578) );
  NAND2_X2 U8417 ( .A1(net247002), .A2(a[11]), .ZN(n6577) );
  AOI21_X2 U8418 ( .B1(n4552), .B2(n6580), .A(n6579), .ZN(n6581) );
  NAND4_X2 U8419 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .ZN(out[11]) );
  INV_X4 U8420 ( .A(n6585), .ZN(n6587) );
  NAND2_X2 U8421 ( .A1(b[12]), .A2(net246788), .ZN(net243374) );
  NAND2_X2 U8422 ( .A1(n6592), .A2(n6591), .ZN(n6887) );
  NAND2_X2 U8423 ( .A1(n6594), .A2(n6593), .ZN(n6883) );
  NAND2_X2 U8424 ( .A1(net246760), .A2(b[16]), .ZN(n6599) );
  INV_X4 U8425 ( .A(n6599), .ZN(n6882) );
  NAND2_X2 U8426 ( .A1(net243774), .A2(net243771), .ZN(n6597) );
  INV_X4 U8427 ( .A(net243771), .ZN(net243769) );
  INV_X4 U8428 ( .A(n6881), .ZN(n6600) );
  INV_X4 U8429 ( .A(net243754), .ZN(net243759) );
  NAND2_X2 U8430 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  INV_X4 U8431 ( .A(n6604), .ZN(n6864) );
  NAND2_X2 U8432 ( .A1(b[17]), .A2(a[24]), .ZN(n6870) );
  NAND2_X2 U8433 ( .A1(a[23]), .A2(b[18]), .ZN(n6606) );
  INV_X4 U8434 ( .A(n6606), .ZN(n6727) );
  NAND2_X2 U8435 ( .A1(net243743), .A2(net243578), .ZN(n6605) );
  OAI21_X2 U8436 ( .B1(net243740), .B2(net243741), .A(n6605), .ZN(n6607) );
  OAI21_X4 U8437 ( .B1(n6608), .B2(n6607), .A(n6606), .ZN(n6861) );
  OAI21_X4 U8438 ( .B1(n4379), .B2(n6729), .A(n6861), .ZN(n6609) );
  XNOR2_X2 U8439 ( .A(n6870), .B(n6609), .ZN(n6877) );
  NAND2_X2 U8440 ( .A1(n6610), .A2(net243731), .ZN(n6611) );
  INV_X4 U8441 ( .A(n6612), .ZN(n6615) );
  OAI21_X4 U8442 ( .B1(n6615), .B2(n6614), .A(n6613), .ZN(n6812) );
  NAND2_X2 U8443 ( .A1(a[14]), .A2(b[27]), .ZN(n6785) );
  INV_X4 U8444 ( .A(n6616), .ZN(n6619) );
  OAI21_X4 U8445 ( .B1(n6619), .B2(n6618), .A(n6617), .ZN(n6783) );
  INV_X4 U8446 ( .A(n6620), .ZN(n6623) );
  OAI21_X4 U8447 ( .B1(n6623), .B2(n6622), .A(n6621), .ZN(n6771) );
  NAND2_X2 U8448 ( .A1(a[10]), .A2(net249231), .ZN(n6971) );
  INV_X4 U8449 ( .A(n6624), .ZN(n6626) );
  NAND2_X2 U8450 ( .A1(n6626), .A2(n6625), .ZN(n6627) );
  OAI21_X4 U8451 ( .B1(n6629), .B2(n6628), .A(n6627), .ZN(n6758) );
  XNOR2_X2 U8452 ( .A(n6971), .B(n6758), .ZN(n6631) );
  NAND2_X2 U8453 ( .A1(a[11]), .A2(net248517), .ZN(n6759) );
  INV_X4 U8454 ( .A(n6759), .ZN(n6630) );
  XNOR2_X2 U8455 ( .A(n6631), .B(n6630), .ZN(n6768) );
  INV_X4 U8456 ( .A(n6768), .ZN(n6642) );
  NAND2_X2 U8457 ( .A1(a[12]), .A2(b[29]), .ZN(n6639) );
  INV_X4 U8458 ( .A(n6639), .ZN(n6637) );
  NAND2_X2 U8459 ( .A1(n6633), .A2(n6632), .ZN(n6634) );
  OAI21_X4 U8460 ( .B1(n6636), .B2(n6635), .A(n6634), .ZN(n6638) );
  NAND2_X2 U8461 ( .A1(n6637), .A2(n6638), .ZN(n6767) );
  INV_X4 U8462 ( .A(n6638), .ZN(n6640) );
  NAND2_X2 U8463 ( .A1(n6767), .A2(n6766), .ZN(n6641) );
  XNOR2_X2 U8464 ( .A(n6642), .B(n6641), .ZN(n6772) );
  NAND2_X2 U8465 ( .A1(a[13]), .A2(net246880), .ZN(n6774) );
  XNOR2_X2 U8466 ( .A(n6772), .B(n6774), .ZN(n6643) );
  XNOR2_X2 U8467 ( .A(n6643), .B(n6771), .ZN(n6781) );
  XNOR2_X2 U8468 ( .A(n6783), .B(n6781), .ZN(n6644) );
  XNOR2_X2 U8469 ( .A(n6644), .B(n6785), .ZN(n6793) );
  INV_X4 U8470 ( .A(n6645), .ZN(n6648) );
  OAI21_X4 U8471 ( .B1(n6648), .B2(n6647), .A(n6646), .ZN(n6792) );
  NAND2_X2 U8472 ( .A1(a[15]), .A2(b[26]), .ZN(n6795) );
  INV_X4 U8473 ( .A(n6649), .ZN(n6652) );
  OAI21_X4 U8474 ( .B1(n6652), .B2(n6651), .A(n6650), .ZN(n6803) );
  NAND2_X2 U8475 ( .A1(a[16]), .A2(b[25]), .ZN(n6805) );
  XNOR2_X2 U8476 ( .A(n6653), .B(n6805), .ZN(n6813) );
  NAND2_X2 U8477 ( .A1(a[17]), .A2(b[24]), .ZN(n6815) );
  XNOR2_X2 U8478 ( .A(n6813), .B(n6815), .ZN(n6654) );
  XNOR2_X2 U8479 ( .A(n6812), .B(n6654), .ZN(n6822) );
  INV_X4 U8480 ( .A(n6655), .ZN(n6658) );
  OAI21_X4 U8481 ( .B1(n6658), .B2(n6657), .A(n6656), .ZN(n6823) );
  XNOR2_X2 U8482 ( .A(n6659), .B(n6823), .ZN(n6836) );
  XNOR2_X2 U8483 ( .A(n4014), .B(n6833), .ZN(n6664) );
  OAI21_X4 U8484 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(n6835) );
  XNOR2_X2 U8485 ( .A(n6664), .B(n6835), .ZN(n6755) );
  INV_X4 U8486 ( .A(n6747), .ZN(n6669) );
  INV_X4 U8487 ( .A(n6665), .ZN(n6668) );
  INV_X4 U8488 ( .A(n6666), .ZN(n6667) );
  OAI21_X4 U8489 ( .B1(n6670), .B2(n6669), .A(n6748), .ZN(n6733) );
  NAND2_X2 U8490 ( .A1(net246836), .A2(a[20]), .ZN(n6754) );
  NAND2_X2 U8491 ( .A1(a[21]), .A2(b[20]), .ZN(n6739) );
  XNOR2_X2 U8492 ( .A(n6754), .B(n6739), .ZN(n6671) );
  FA_X1 U8493 ( .A(n6671), .B(n6733), .CI(n6755), .S(n6676) );
  NAND2_X2 U8494 ( .A1(n6674), .A2(n6672), .ZN(n6737) );
  NAND2_X2 U8495 ( .A1(n6673), .A2(n6672), .ZN(n6736) );
  NAND2_X2 U8496 ( .A1(n6674), .A2(n6673), .ZN(n6738) );
  XNOR2_X2 U8497 ( .A(n6676), .B(n6675), .ZN(n6851) );
  NAND2_X2 U8498 ( .A1(b[19]), .A2(a[22]), .ZN(n6848) );
  XNOR2_X2 U8499 ( .A(n6851), .B(n6848), .ZN(n6677) );
  XNOR2_X2 U8500 ( .A(n6850), .B(n6677), .ZN(n6876) );
  XNOR2_X2 U8501 ( .A(n4402), .B(n6878), .ZN(net243403) );
  XNOR2_X2 U8502 ( .A(net248444), .B(net243634), .ZN(n6893) );
  NAND2_X2 U8503 ( .A1(b[13]), .A2(a[28]), .ZN(n6888) );
  XNOR2_X2 U8504 ( .A(n6893), .B(n6888), .ZN(n6685) );
  XNOR2_X2 U8505 ( .A(n6685), .B(n6686), .ZN(net243371) );
  INV_X4 U8506 ( .A(n6687), .ZN(n6688) );
  NOR3_X4 U8507 ( .A1(n6688), .A2(net246812), .A3(net243628), .ZN(net243367)
         );
  NAND2_X2 U8508 ( .A1(b[11]), .A2(a[30]), .ZN(net243368) );
  XNOR2_X2 U8509 ( .A(net243367), .B(net243368), .ZN(n6689) );
  XNOR2_X2 U8510 ( .A(net243625), .B(n6689), .ZN(n6692) );
  NAND2_X2 U8511 ( .A1(net240913), .A2(net243587), .ZN(n6691) );
  NAND2_X2 U8512 ( .A1(n6691), .A2(n4550), .ZN(n6710) );
  INV_X4 U8513 ( .A(n6693), .ZN(n6694) );
  AOI21_X4 U8514 ( .B1(n4557), .B2(n7415), .A(n3992), .ZN(n6698) );
  OAI221_X2 U8515 ( .B1(n1386), .B2(n4533), .C1(n853), .C2(n8115), .A(n6698), 
        .ZN(n6908) );
  NAND2_X2 U8516 ( .A1(n4558), .A2(n7039), .ZN(n6704) );
  NAND2_X2 U8517 ( .A1(n6699), .A2(n6564), .ZN(n6703) );
  NAND2_X2 U8518 ( .A1(n4554), .A2(n7419), .ZN(n6702) );
  NAND2_X2 U8519 ( .A1(n7825), .A2(n4565), .ZN(n6701) );
  NAND4_X2 U8520 ( .A1(n6704), .A2(n6703), .A3(n6702), .A4(n6701), .ZN(n6909)
         );
  INV_X4 U8521 ( .A(n6909), .ZN(n6705) );
  AOI21_X2 U8522 ( .B1(n8125), .B2(n6908), .A(n6706), .ZN(n6707) );
  XNOR2_X2 U8523 ( .A(net246926), .B(b[10]), .ZN(n6902) );
  XNOR2_X2 U8524 ( .A(a[10]), .B(n6902), .ZN(n6717) );
  INV_X4 U8525 ( .A(n6711), .ZN(n6715) );
  NAND2_X2 U8526 ( .A1(n6713), .A2(n6712), .ZN(n6714) );
  OAI21_X4 U8527 ( .B1(n6716), .B2(n6715), .A(n6714), .ZN(n6903) );
  XNOR2_X2 U8528 ( .A(n6717), .B(n6903), .ZN(n6721) );
  NAND2_X2 U8529 ( .A1(n8784), .A2(n6718), .ZN(n6719) );
  AOI21_X2 U8530 ( .B1(n4552), .B2(n6721), .A(n6720), .ZN(n6722) );
  OAI211_X2 U8531 ( .C1(n6724), .C2(net243587), .A(n6723), .B(n6722), .ZN(
        out[10]) );
  NAND3_X4 U8532 ( .A1(b[10]), .A2(a[31]), .A3(n6725), .ZN(n7018) );
  NAND2_X2 U8533 ( .A1(b[10]), .A2(a[30]), .ZN(n7017) );
  XNOR2_X2 U8534 ( .A(n7015), .B(n7017), .ZN(n6895) );
  INV_X4 U8535 ( .A(n6729), .ZN(n6731) );
  NAND2_X2 U8536 ( .A1(a[22]), .A2(b[18]), .ZN(n6944) );
  XNOR2_X2 U8537 ( .A(n6946), .B(n6944), .ZN(net243439) );
  XNOR2_X2 U8538 ( .A(n6735), .B(n6734), .ZN(n6741) );
  NAND3_X2 U8539 ( .A1(n6738), .A2(n6737), .A3(n6736), .ZN(n6740) );
  NAND2_X2 U8540 ( .A1(n6741), .A2(n6740), .ZN(n6743) );
  XNOR2_X2 U8541 ( .A(n6957), .B(n7089), .ZN(n6847) );
  INV_X4 U8542 ( .A(n6754), .ZN(n6752) );
  XNOR2_X2 U8543 ( .A(n6744), .B(n6833), .ZN(n6745) );
  XNOR2_X2 U8544 ( .A(n6745), .B(n6835), .ZN(n6751) );
  NAND2_X2 U8545 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  NAND2_X2 U8546 ( .A1(a[19]), .A2(net246836), .ZN(n6959) );
  INV_X4 U8547 ( .A(n6959), .ZN(n6757) );
  OAI22_X2 U8548 ( .A1(n6960), .A2(n6959), .B1(n6756), .B2(n6757), .ZN(n6845)
         );
  NAND2_X2 U8549 ( .A1(a[11]), .A2(b[29]), .ZN(n6976) );
  INV_X4 U8550 ( .A(n6969), .ZN(n6765) );
  INV_X4 U8551 ( .A(n6758), .ZN(n6760) );
  NAND2_X2 U8552 ( .A1(n6760), .A2(n6759), .ZN(n6762) );
  OAI21_X4 U8553 ( .B1(n6760), .B2(n6759), .A(n6971), .ZN(n6761) );
  NAND2_X2 U8554 ( .A1(n6762), .A2(n6761), .ZN(n6970) );
  INV_X4 U8555 ( .A(n6970), .ZN(n6763) );
  NAND2_X2 U8556 ( .A1(n6763), .A2(n3958), .ZN(n6968) );
  OAI21_X4 U8557 ( .B1(n6763), .B2(n3958), .A(n6968), .ZN(n6764) );
  XNOR2_X2 U8558 ( .A(n6765), .B(n6764), .ZN(n6973) );
  INV_X4 U8559 ( .A(n6766), .ZN(n6769) );
  OAI21_X4 U8560 ( .B1(n6769), .B2(n6768), .A(n6767), .ZN(n6974) );
  XNOR2_X2 U8561 ( .A(n6973), .B(n6974), .ZN(n6770) );
  XNOR2_X2 U8562 ( .A(n6976), .B(n6770), .ZN(n6966) );
  NAND2_X2 U8563 ( .A1(a[12]), .A2(net246880), .ZN(n6778) );
  INV_X4 U8564 ( .A(n6778), .ZN(n6776) );
  NAND2_X2 U8565 ( .A1(n4388), .A2(n6771), .ZN(n6773) );
  OAI21_X4 U8566 ( .B1(n6775), .B2(n6774), .A(n6773), .ZN(n6777) );
  NAND2_X2 U8567 ( .A1(n6776), .A2(n6777), .ZN(n6965) );
  INV_X4 U8568 ( .A(n6777), .ZN(n6779) );
  NAND2_X2 U8569 ( .A1(n6779), .A2(n6778), .ZN(n6964) );
  NAND2_X2 U8570 ( .A1(n6965), .A2(n6964), .ZN(n6780) );
  XNOR2_X2 U8571 ( .A(n6966), .B(n6780), .ZN(n6983) );
  NAND2_X2 U8572 ( .A1(a[13]), .A2(b[27]), .ZN(n6789) );
  INV_X4 U8573 ( .A(n6789), .ZN(n6787) );
  INV_X4 U8574 ( .A(n6781), .ZN(n6782) );
  OAI21_X4 U8575 ( .B1(n6786), .B2(n6785), .A(n6784), .ZN(n6788) );
  NAND2_X2 U8576 ( .A1(n6787), .A2(n6788), .ZN(n6982) );
  INV_X4 U8577 ( .A(n6788), .ZN(n6790) );
  NAND2_X2 U8578 ( .A1(n6790), .A2(n6789), .ZN(n6981) );
  XNOR2_X2 U8579 ( .A(n6983), .B(n6791), .ZN(n6987) );
  NAND2_X2 U8580 ( .A1(a[14]), .A2(b[26]), .ZN(n6799) );
  INV_X4 U8581 ( .A(n6799), .ZN(n6797) );
  NAND2_X2 U8582 ( .A1(n6797), .A2(n6798), .ZN(n6986) );
  INV_X4 U8583 ( .A(n6798), .ZN(n6800) );
  XNOR2_X2 U8584 ( .A(n6987), .B(n6801), .ZN(n6991) );
  NAND2_X2 U8585 ( .A1(a[15]), .A2(b[25]), .ZN(n6809) );
  INV_X4 U8586 ( .A(n6809), .ZN(n6807) );
  NAND2_X2 U8587 ( .A1(n6807), .A2(n6808), .ZN(n6990) );
  INV_X4 U8588 ( .A(n6808), .ZN(n6810) );
  NAND2_X2 U8589 ( .A1(n6990), .A2(n6989), .ZN(n6811) );
  XNOR2_X2 U8590 ( .A(n6991), .B(n6811), .ZN(n6995) );
  NAND2_X2 U8591 ( .A1(a[16]), .A2(b[24]), .ZN(n6819) );
  INV_X4 U8592 ( .A(n6819), .ZN(n6817) );
  OAI21_X4 U8593 ( .B1(n6816), .B2(n6815), .A(n6814), .ZN(n6818) );
  NAND2_X2 U8594 ( .A1(n6817), .A2(n6818), .ZN(n6994) );
  INV_X4 U8595 ( .A(n6818), .ZN(n6820) );
  NAND2_X2 U8596 ( .A1(n6820), .A2(n6819), .ZN(n6993) );
  NAND2_X2 U8597 ( .A1(n6994), .A2(n6993), .ZN(n6821) );
  XNOR2_X2 U8598 ( .A(n6995), .B(n6821), .ZN(n7000) );
  NAND2_X2 U8599 ( .A1(a[17]), .A2(b[23]), .ZN(n6830) );
  INV_X4 U8600 ( .A(n6830), .ZN(n6828) );
  NAND2_X2 U8601 ( .A1(n6824), .A2(n6823), .ZN(n6825) );
  OAI21_X4 U8602 ( .B1(n6827), .B2(n6826), .A(n6825), .ZN(n6829) );
  NAND2_X2 U8603 ( .A1(n6828), .A2(n6829), .ZN(n6999) );
  INV_X4 U8604 ( .A(n6829), .ZN(n6831) );
  NAND2_X2 U8605 ( .A1(n6831), .A2(n6830), .ZN(n6998) );
  NAND2_X2 U8606 ( .A1(n6999), .A2(n6998), .ZN(n6832) );
  XNOR2_X2 U8607 ( .A(n7000), .B(n6832), .ZN(n7005) );
  INV_X4 U8608 ( .A(n7005), .ZN(n6844) );
  INV_X4 U8609 ( .A(n6841), .ZN(n6839) );
  INV_X4 U8610 ( .A(n6833), .ZN(n6834) );
  NAND2_X2 U8611 ( .A1(a[18]), .A2(b[22]), .ZN(n6842) );
  INV_X4 U8612 ( .A(n6842), .ZN(n6837) );
  OAI21_X4 U8613 ( .B1(n6839), .B2(n6838), .A(n6837), .ZN(n7004) );
  XNOR2_X2 U8614 ( .A(n6844), .B(n6843), .ZN(n6962) );
  XNOR2_X2 U8615 ( .A(n6845), .B(n6962), .ZN(n7091) );
  XNOR2_X2 U8616 ( .A(n6847), .B(n6846), .ZN(n6955) );
  INV_X4 U8617 ( .A(n6955), .ZN(n6860) );
  NAND2_X2 U8618 ( .A1(b[19]), .A2(a[21]), .ZN(n6857) );
  INV_X4 U8619 ( .A(n6857), .ZN(n6855) );
  INV_X4 U8620 ( .A(n6848), .ZN(n6849) );
  NAND2_X2 U8621 ( .A1(n6849), .A2(n6850), .ZN(n6853) );
  NAND3_X2 U8622 ( .A1(n6854), .A2(n6853), .A3(n6852), .ZN(n6856) );
  NAND2_X2 U8623 ( .A1(n6855), .A2(n6856), .ZN(n6954) );
  INV_X4 U8624 ( .A(n6856), .ZN(n6858) );
  NAND2_X2 U8625 ( .A1(n6858), .A2(n6857), .ZN(n6953) );
  NAND2_X2 U8626 ( .A1(n6954), .A2(n6953), .ZN(n6859) );
  XNOR2_X2 U8627 ( .A(n6860), .B(n6859), .ZN(net243261) );
  NAND2_X2 U8628 ( .A1(b[17]), .A2(a[23]), .ZN(n6872) );
  INV_X4 U8629 ( .A(n6872), .ZN(n6943) );
  XNOR2_X2 U8630 ( .A(n6863), .B(n6876), .ZN(n6871) );
  INV_X4 U8631 ( .A(n6870), .ZN(n6867) );
  NAND2_X2 U8632 ( .A1(n6867), .A2(n6866), .ZN(n6868) );
  INV_X4 U8633 ( .A(n6942), .ZN(n6873) );
  INV_X4 U8634 ( .A(net243423), .ZN(net243422) );
  NOR2_X4 U8635 ( .A1(n6882), .A2(net243422), .ZN(n6875) );
  XNOR2_X2 U8636 ( .A(n6678), .B(n6878), .ZN(n6879) );
  NAND2_X2 U8637 ( .A1(b[15]), .A2(net246760), .ZN(net243291) );
  INV_X4 U8638 ( .A(net243395), .ZN(net243398) );
  NAND2_X2 U8639 ( .A1(n6887), .A2(n6888), .ZN(n6886) );
  INV_X4 U8640 ( .A(n6887), .ZN(n6891) );
  INV_X4 U8641 ( .A(n6888), .ZN(n6889) );
  NAND2_X2 U8642 ( .A1(b[13]), .A2(net246772), .ZN(net243310) );
  XNOR2_X2 U8643 ( .A(n6895), .B(net242899), .ZN(n6935) );
  NAND2_X2 U8644 ( .A1(net240782), .A2(a[9]), .ZN(n6896) );
  NAND2_X2 U8645 ( .A1(b[9]), .A2(n6897), .ZN(n6934) );
  NAND2_X2 U8646 ( .A1(net240913), .A2(net243356), .ZN(n6898) );
  NAND2_X2 U8647 ( .A1(n6898), .A2(n4550), .ZN(n6899) );
  NAND2_X2 U8648 ( .A1(n8784), .A2(n6900), .ZN(n6932) );
  NAND2_X2 U8649 ( .A1(n6903), .A2(n6901), .ZN(n6906) );
  INV_X4 U8650 ( .A(n6902), .ZN(n6905) );
  INV_X4 U8651 ( .A(n6903), .ZN(n6904) );
  AOI22_X2 U8652 ( .A1(n6906), .A2(n6905), .B1(n6904), .B2(a[10]), .ZN(n7030)
         );
  XNOR2_X2 U8653 ( .A(net246924), .B(b[9]), .ZN(n7028) );
  XNOR2_X2 U8654 ( .A(a[9]), .B(n7028), .ZN(n6907) );
  XNOR2_X2 U8655 ( .A(n7030), .B(n6907), .ZN(n6930) );
  INV_X4 U8656 ( .A(n6908), .ZN(n6911) );
  NAND2_X2 U8657 ( .A1(n8841), .A2(n6909), .ZN(n6910) );
  INV_X4 U8658 ( .A(n8300), .ZN(n6912) );
  NAND2_X2 U8659 ( .A1(n7044), .A2(n6912), .ZN(n8111) );
  INV_X4 U8660 ( .A(n8111), .ZN(n6915) );
  OAI221_X2 U8661 ( .B1(n6915), .B2(n4533), .C1(n949), .C2(n8832), .A(n6914), 
        .ZN(n6916) );
  INV_X4 U8662 ( .A(n6916), .ZN(n7047) );
  NAND2_X2 U8663 ( .A1(net247082), .A2(net246760), .ZN(n6917) );
  NAND2_X2 U8664 ( .A1(n8118), .A2(n4565), .ZN(n6923) );
  NAND2_X2 U8665 ( .A1(n4554), .A2(n7658), .ZN(n6922) );
  AOI22_X2 U8666 ( .A1(n4561), .A2(n6920), .B1(n4557), .B2(n7247), .ZN(n6921)
         );
  NAND3_X2 U8667 ( .A1(n6923), .A2(n6922), .A3(n6921), .ZN(n7035) );
  NAND2_X2 U8668 ( .A1(n8318), .A2(n7035), .ZN(n6924) );
  NOR2_X4 U8669 ( .A1(n6926), .A2(n6925), .ZN(n6928) );
  NAND2_X2 U8670 ( .A1(net247002), .A2(a[9]), .ZN(n6927) );
  AOI21_X2 U8671 ( .B1(n4552), .B2(n6930), .A(n6929), .ZN(n6931) );
  NAND4_X2 U8672 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(out[9])
         );
  INV_X4 U8673 ( .A(n7232), .ZN(n7229) );
  NAND2_X2 U8674 ( .A1(b[9]), .A2(a[30]), .ZN(n7231) );
  XNOR2_X2 U8675 ( .A(n7229), .B(n7231), .ZN(net243159) );
  NAND2_X2 U8676 ( .A1(b[13]), .A2(net246766), .ZN(n7224) );
  INV_X4 U8677 ( .A(n7224), .ZN(n7227) );
  NOR2_X4 U8678 ( .A1(net243298), .A2(net243299), .ZN(net243296) );
  INV_X4 U8679 ( .A(net243292), .ZN(net243289) );
  NAND2_X2 U8680 ( .A1(net243283), .A2(net243284), .ZN(n6937) );
  OAI21_X4 U8681 ( .B1(n6938), .B2(net243281), .A(n6937), .ZN(n7217) );
  INV_X4 U8682 ( .A(n7221), .ZN(n7218) );
  OAI22_X2 U8683 ( .A1(n7222), .A2(n7221), .B1(n7218), .B2(n7217), .ZN(n7014)
         );
  NAND2_X2 U8684 ( .A1(b[15]), .A2(net246754), .ZN(net243081) );
  XNOR2_X2 U8685 ( .A(net243278), .B(net243081), .ZN(n7013) );
  INV_X4 U8686 ( .A(net243270), .ZN(net243268) );
  NAND2_X2 U8687 ( .A1(n6941), .A2(n7072), .ZN(n7371) );
  NAND2_X2 U8688 ( .A1(b[17]), .A2(a[22]), .ZN(n7078) );
  NAND2_X2 U8689 ( .A1(a[21]), .A2(b[18]), .ZN(n6949) );
  INV_X4 U8690 ( .A(n6949), .ZN(n6948) );
  INV_X4 U8691 ( .A(n6944), .ZN(n6945) );
  NAND2_X2 U8692 ( .A1(n6945), .A2(net243261), .ZN(n6951) );
  NAND2_X2 U8693 ( .A1(n4417), .A2(net243261), .ZN(n6952) );
  NAND4_X2 U8694 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(n6949), .ZN(n7085)
         );
  INV_X4 U8695 ( .A(n6953), .ZN(n6956) );
  OAI21_X4 U8696 ( .B1(n6956), .B2(n6955), .A(n6954), .ZN(n7208) );
  NAND2_X2 U8697 ( .A1(b[19]), .A2(a[20]), .ZN(n7206) );
  XNOR2_X2 U8698 ( .A(n7208), .B(n7206), .ZN(n7084) );
  INV_X4 U8699 ( .A(n6957), .ZN(n7090) );
  NAND2_X2 U8700 ( .A1(a[18]), .A2(net246836), .ZN(n7197) );
  NAND2_X2 U8701 ( .A1(n6960), .A2(n6959), .ZN(n6961) );
  OAI21_X4 U8702 ( .B1(n6963), .B2(n6962), .A(n6961), .ZN(n7194) );
  XNOR2_X2 U8703 ( .A(n7197), .B(n7194), .ZN(n7008) );
  INV_X4 U8704 ( .A(n6964), .ZN(n6967) );
  OAI21_X4 U8705 ( .B1(n6967), .B2(n6966), .A(n6965), .ZN(n7124) );
  NAND2_X2 U8706 ( .A1(a[9]), .A2(net246902), .ZN(n7105) );
  OAI221_X2 U8707 ( .B1(n7105), .B2(n6971), .C1(n6970), .C2(n6969), .A(n6968), 
        .ZN(n7104) );
  NAND2_X2 U8708 ( .A1(a[8]), .A2(net246916), .ZN(n7318) );
  XNOR2_X2 U8709 ( .A(n7105), .B(n7318), .ZN(n6972) );
  XNOR2_X2 U8710 ( .A(n7104), .B(n6972), .ZN(n7114) );
  NAND2_X2 U8711 ( .A1(n6974), .A2(n6973), .ZN(n6975) );
  OAI21_X4 U8712 ( .B1(n6977), .B2(n6976), .A(n6975), .ZN(n7115) );
  XOR2_X2 U8713 ( .A(n7114), .B(n7115), .Z(n6978) );
  NAND2_X2 U8714 ( .A1(a[10]), .A2(b[29]), .ZN(n7117) );
  XNOR2_X2 U8715 ( .A(n6978), .B(n7117), .ZN(n7125) );
  NAND2_X2 U8716 ( .A1(a[11]), .A2(net246880), .ZN(n7127) );
  INV_X4 U8717 ( .A(n7127), .ZN(n6979) );
  XNOR2_X2 U8718 ( .A(n7125), .B(n6979), .ZN(n6980) );
  XNOR2_X2 U8719 ( .A(n7124), .B(n6980), .ZN(n7135) );
  INV_X4 U8720 ( .A(n6981), .ZN(n6984) );
  OAI21_X4 U8721 ( .B1(n6984), .B2(n6983), .A(n6982), .ZN(n7134) );
  NAND2_X2 U8722 ( .A1(a[12]), .A2(b[27]), .ZN(n7137) );
  INV_X4 U8723 ( .A(n6985), .ZN(n6988) );
  OAI21_X4 U8724 ( .B1(n6988), .B2(n6987), .A(n6986), .ZN(n7144) );
  NAND2_X2 U8725 ( .A1(a[13]), .A2(b[26]), .ZN(n7147) );
  INV_X4 U8726 ( .A(n6989), .ZN(n6992) );
  OAI21_X4 U8727 ( .B1(n6992), .B2(n6991), .A(n6990), .ZN(n7155) );
  NAND2_X2 U8728 ( .A1(a[14]), .A2(b[25]), .ZN(n7157) );
  NAND2_X2 U8729 ( .A1(a[15]), .A2(b[24]), .ZN(n7167) );
  INV_X4 U8730 ( .A(n6993), .ZN(n6996) );
  OAI21_X4 U8731 ( .B1(n6996), .B2(n6995), .A(n6994), .ZN(n7164) );
  XNOR2_X2 U8732 ( .A(n6997), .B(n7164), .ZN(n7175) );
  NAND2_X2 U8733 ( .A1(a[16]), .A2(b[23]), .ZN(n7177) );
  INV_X4 U8734 ( .A(n6998), .ZN(n7001) );
  OAI21_X4 U8735 ( .B1(n7001), .B2(n7000), .A(n6999), .ZN(n7174) );
  XNOR2_X2 U8736 ( .A(n7002), .B(n7174), .ZN(n7185) );
  NAND2_X2 U8737 ( .A1(a[17]), .A2(b[22]), .ZN(n7187) );
  XNOR2_X2 U8738 ( .A(n7185), .B(n7187), .ZN(n7007) );
  INV_X4 U8739 ( .A(n7003), .ZN(n7006) );
  XNOR2_X2 U8740 ( .A(n7008), .B(n4455), .ZN(n7097) );
  NAND2_X2 U8741 ( .A1(a[19]), .A2(b[20]), .ZN(n7100) );
  XNOR2_X2 U8742 ( .A(n7097), .B(n7100), .ZN(n7009) );
  XNOR2_X2 U8743 ( .A(n7098), .B(n7009), .ZN(n7205) );
  XNOR2_X2 U8744 ( .A(n7084), .B(n7205), .ZN(n7076) );
  XNOR2_X2 U8745 ( .A(n7010), .B(n7082), .ZN(n7372) );
  XNOR2_X2 U8746 ( .A(n7011), .B(n7372), .ZN(n7012) );
  XNOR2_X2 U8747 ( .A(n7013), .B(n7012), .ZN(n7219) );
  XNOR2_X2 U8748 ( .A(n7219), .B(n7014), .ZN(net242909) );
  INV_X4 U8749 ( .A(net243184), .ZN(net243182) );
  NAND2_X2 U8750 ( .A1(b[12]), .A2(net246772), .ZN(net243119) );
  INV_X4 U8751 ( .A(n7017), .ZN(n7016) );
  NAND2_X2 U8752 ( .A1(n7016), .A2(n7015), .ZN(net242900) );
  INV_X4 U8753 ( .A(net242900), .ZN(net243171) );
  NAND2_X2 U8754 ( .A1(b[10]), .A2(net246788), .ZN(net242894) );
  NAND2_X2 U8755 ( .A1(n7018), .A2(n7017), .ZN(net243166) );
  NAND2_X2 U8756 ( .A1(net243167), .A2(net243168), .ZN(n7020) );
  INV_X4 U8757 ( .A(net243166), .ZN(net242898) );
  NAND3_X2 U8758 ( .A1(n7021), .A2(n7020), .A3(n7019), .ZN(n7022) );
  XNOR2_X2 U8759 ( .A(n7022), .B(net248775), .ZN(net242672) );
  NAND2_X2 U8760 ( .A1(net240782), .A2(a[8]), .ZN(n7023) );
  NAND2_X2 U8761 ( .A1(b[8]), .A2(n7024), .ZN(n7058) );
  NAND2_X2 U8762 ( .A1(net240913), .A2(net242878), .ZN(n7025) );
  NAND2_X2 U8763 ( .A1(n7025), .A2(n4550), .ZN(n7026) );
  NAND2_X2 U8764 ( .A1(n8784), .A2(n7027), .ZN(n7056) );
  XNOR2_X2 U8765 ( .A(net246924), .B(b[8]), .ZN(n7241) );
  XNOR2_X2 U8766 ( .A(a[8]), .B(n7241), .ZN(n7034) );
  INV_X4 U8767 ( .A(n7028), .ZN(n7032) );
  NAND2_X2 U8768 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  OAI21_X4 U8769 ( .B1(n7033), .B2(n7032), .A(n7031), .ZN(n7242) );
  XNOR2_X2 U8770 ( .A(n7034), .B(n7242), .ZN(n7054) );
  INV_X4 U8771 ( .A(n7035), .ZN(n7043) );
  NAND2_X2 U8772 ( .A1(net247082), .A2(net246754), .ZN(n7036) );
  NAND3_X2 U8773 ( .A1(n7038), .A2(n7037), .A3(n7036), .ZN(n8305) );
  NAND2_X2 U8774 ( .A1(n8305), .A2(n4565), .ZN(n7042) );
  NAND2_X2 U8775 ( .A1(n4554), .A2(n7825), .ZN(n7041) );
  AOI22_X2 U8776 ( .A1(n4561), .A2(n7039), .B1(n4557), .B2(n7419), .ZN(n7040)
         );
  OAI22_X2 U8777 ( .A1(n7043), .A2(n4539), .B1(n3984), .B2(n4537), .ZN(n7050)
         );
  OAI21_X4 U8778 ( .B1(net246956), .B2(net240852), .A(n7044), .ZN(n8314) );
  AOI22_X2 U8779 ( .A1(n4555), .A2(n7415), .B1(n4561), .B2(n8314), .ZN(n7045)
         );
  OAI221_X2 U8780 ( .B1(n1386), .B2(n8832), .C1(n853), .C2(n4566), .A(n7045), 
        .ZN(n7046) );
  INV_X4 U8781 ( .A(n7046), .ZN(n7255) );
  NOR3_X4 U8782 ( .A1(n7050), .A2(n7049), .A3(n7048), .ZN(n7052) );
  NAND2_X2 U8783 ( .A1(net247002), .A2(a[8]), .ZN(n7051) );
  AOI21_X2 U8784 ( .B1(n4552), .B2(n7054), .A(n7053), .ZN(n7055) );
  NAND4_X2 U8785 ( .A1(n7058), .A2(n7057), .A3(n7056), .A4(n7055), .ZN(out[8])
         );
  NAND2_X2 U8786 ( .A1(b[12]), .A2(net246766), .ZN(net242824) );
  INV_X4 U8787 ( .A(net243099), .ZN(net243079) );
  NOR2_X2 U8788 ( .A1(net243079), .A2(net243098), .ZN(n7071) );
  XNOR2_X2 U8789 ( .A(net243093), .B(n7077), .ZN(n7061) );
  INV_X4 U8790 ( .A(n7076), .ZN(n7059) );
  INV_X4 U8791 ( .A(n7078), .ZN(n7080) );
  INV_X4 U8792 ( .A(n7062), .ZN(n7066) );
  AOI21_X2 U8793 ( .B1(n7064), .B2(n7063), .A(n7073), .ZN(n7065) );
  NOR2_X4 U8794 ( .A1(n7066), .A2(n7065), .ZN(n7067) );
  XNOR2_X2 U8795 ( .A(n7068), .B(n7067), .ZN(n7070) );
  INV_X4 U8796 ( .A(net243081), .ZN(net243080) );
  OAI21_X4 U8797 ( .B1(net243078), .B2(net243079), .A(net243080), .ZN(n7069)
         );
  OAI21_X4 U8798 ( .B1(n7071), .B2(n7070), .A(n7069), .ZN(n7286) );
  INV_X4 U8799 ( .A(n7286), .ZN(n7283) );
  NAND2_X2 U8800 ( .A1(b[15]), .A2(a[23]), .ZN(n7282) );
  INV_X4 U8801 ( .A(n7282), .ZN(n7287) );
  NAND2_X2 U8802 ( .A1(a[22]), .A2(b[16]), .ZN(n7374) );
  XNOR2_X2 U8803 ( .A(n7075), .B(n7374), .ZN(n7214) );
  XNOR2_X2 U8804 ( .A(n7077), .B(n7076), .ZN(n7082) );
  INV_X4 U8805 ( .A(n7361), .ZN(n7081) );
  AOI21_X4 U8806 ( .B1(n7082), .B2(n7359), .A(n7081), .ZN(n7364) );
  NAND2_X2 U8807 ( .A1(b[17]), .A2(a[21]), .ZN(n7363) );
  OAI21_X2 U8808 ( .B1(n7364), .B2(n7363), .A(n7083), .ZN(n7213) );
  XNOR2_X2 U8809 ( .A(n7205), .B(n7084), .ZN(n7086) );
  NAND2_X2 U8810 ( .A1(n7086), .A2(n7085), .ZN(n7088) );
  NAND2_X2 U8811 ( .A1(a[20]), .A2(b[18]), .ZN(n7292) );
  XNOR2_X2 U8812 ( .A(n7289), .B(n7292), .ZN(n7212) );
  INV_X4 U8813 ( .A(n7089), .ZN(n7092) );
  NAND2_X2 U8814 ( .A1(n7090), .A2(n7092), .ZN(n7095) );
  NAND2_X2 U8815 ( .A1(n7092), .A2(n7091), .ZN(n7093) );
  NAND3_X2 U8816 ( .A1(n7095), .A2(n7094), .A3(n7093), .ZN(n7096) );
  NAND2_X2 U8817 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  OAI21_X4 U8818 ( .B1(n7101), .B2(n7100), .A(n7099), .ZN(n7301) );
  NAND2_X2 U8819 ( .A1(a[18]), .A2(b[20]), .ZN(n7102) );
  INV_X4 U8820 ( .A(n7102), .ZN(n7302) );
  OAI22_X2 U8821 ( .A1(n7103), .A2(n7102), .B1(n7302), .B2(n7301), .ZN(n7204)
         );
  INV_X4 U8822 ( .A(n7104), .ZN(n7106) );
  NAND2_X2 U8823 ( .A1(n7106), .A2(n7105), .ZN(n7108) );
  OAI21_X4 U8824 ( .B1(n7106), .B2(n7105), .A(n7318), .ZN(n7107) );
  NAND2_X2 U8825 ( .A1(n7108), .A2(n7107), .ZN(n7110) );
  INV_X4 U8826 ( .A(n7110), .ZN(n7316) );
  NAND2_X2 U8827 ( .A1(a[8]), .A2(net248517), .ZN(n7111) );
  INV_X4 U8828 ( .A(n7111), .ZN(n7109) );
  NAND2_X2 U8829 ( .A1(n7316), .A2(n7109), .ZN(n7319) );
  NAND2_X2 U8830 ( .A1(n7111), .A2(n7110), .ZN(n7112) );
  NAND2_X2 U8831 ( .A1(n7319), .A2(n7112), .ZN(n7113) );
  XNOR2_X2 U8832 ( .A(n7315), .B(n7113), .ZN(n7324) );
  NAND2_X2 U8833 ( .A1(a[9]), .A2(b[29]), .ZN(n7121) );
  INV_X4 U8834 ( .A(n7121), .ZN(n7119) );
  OAI21_X4 U8835 ( .B1(n7118), .B2(n7117), .A(n7116), .ZN(n7120) );
  INV_X4 U8836 ( .A(n7120), .ZN(n7122) );
  NAND2_X2 U8837 ( .A1(n7122), .A2(n7121), .ZN(n7322) );
  NAND2_X2 U8838 ( .A1(n7323), .A2(n7322), .ZN(n7123) );
  XNOR2_X2 U8839 ( .A(n7324), .B(n7123), .ZN(n7329) );
  NAND2_X2 U8840 ( .A1(a[10]), .A2(net246880), .ZN(n7131) );
  INV_X4 U8841 ( .A(n7131), .ZN(n7129) );
  INV_X4 U8842 ( .A(n7130), .ZN(n7132) );
  XNOR2_X2 U8843 ( .A(n7329), .B(n7133), .ZN(n7333) );
  NAND2_X2 U8844 ( .A1(a[11]), .A2(b[27]), .ZN(n7141) );
  INV_X4 U8845 ( .A(n7141), .ZN(n7139) );
  OAI21_X4 U8846 ( .B1(n7138), .B2(n7137), .A(n7136), .ZN(n7140) );
  NAND2_X2 U8847 ( .A1(n7139), .A2(n7140), .ZN(n7332) );
  INV_X4 U8848 ( .A(n7140), .ZN(n7142) );
  NAND2_X2 U8849 ( .A1(n7142), .A2(n7141), .ZN(n7331) );
  NAND2_X2 U8850 ( .A1(n7332), .A2(n7331), .ZN(n7143) );
  XNOR2_X2 U8851 ( .A(n7333), .B(n7143), .ZN(n7337) );
  NAND2_X2 U8852 ( .A1(a[12]), .A2(b[26]), .ZN(n7151) );
  INV_X4 U8853 ( .A(n7151), .ZN(n7149) );
  NAND2_X2 U8854 ( .A1(n7149), .A2(n7150), .ZN(n7336) );
  INV_X4 U8855 ( .A(n7150), .ZN(n7152) );
  NAND2_X2 U8856 ( .A1(n7152), .A2(n7151), .ZN(n7335) );
  NAND2_X2 U8857 ( .A1(n7336), .A2(n7335), .ZN(n7153) );
  XNOR2_X2 U8858 ( .A(n7337), .B(n7153), .ZN(n7342) );
  NAND2_X2 U8859 ( .A1(a[13]), .A2(b[25]), .ZN(n7161) );
  INV_X4 U8860 ( .A(n7161), .ZN(n7159) );
  OAI21_X4 U8861 ( .B1(n7158), .B2(n7157), .A(n7156), .ZN(n7160) );
  NAND2_X2 U8862 ( .A1(n7159), .A2(n7160), .ZN(n7341) );
  INV_X4 U8863 ( .A(n7160), .ZN(n7162) );
  NAND2_X2 U8864 ( .A1(n7162), .A2(n7161), .ZN(n7340) );
  NAND2_X2 U8865 ( .A1(n7341), .A2(n7340), .ZN(n7163) );
  XNOR2_X2 U8866 ( .A(n7342), .B(n7163), .ZN(n7346) );
  NAND2_X2 U8867 ( .A1(a[14]), .A2(b[24]), .ZN(n7171) );
  INV_X4 U8868 ( .A(n7171), .ZN(n7169) );
  OAI21_X4 U8869 ( .B1(n7168), .B2(n7167), .A(n7166), .ZN(n7170) );
  NAND2_X2 U8870 ( .A1(n7169), .A2(n7170), .ZN(n7345) );
  INV_X4 U8871 ( .A(n7170), .ZN(n7172) );
  NAND2_X2 U8872 ( .A1(n7172), .A2(n7171), .ZN(n7344) );
  NAND2_X2 U8873 ( .A1(n7345), .A2(n7344), .ZN(n7173) );
  XNOR2_X2 U8874 ( .A(n7346), .B(n7173), .ZN(n7352) );
  NAND2_X2 U8875 ( .A1(a[15]), .A2(b[23]), .ZN(n7181) );
  INV_X4 U8876 ( .A(n7181), .ZN(n7179) );
  OAI21_X4 U8877 ( .B1(n7178), .B2(n7177), .A(n7176), .ZN(n7180) );
  NAND2_X2 U8878 ( .A1(n7179), .A2(n7180), .ZN(n7351) );
  INV_X4 U8879 ( .A(n7180), .ZN(n7182) );
  NAND2_X2 U8880 ( .A1(n7182), .A2(n7181), .ZN(n7350) );
  NAND2_X2 U8881 ( .A1(n7351), .A2(n7350), .ZN(n7183) );
  XNOR2_X2 U8882 ( .A(n7352), .B(n7183), .ZN(n7313) );
  NAND2_X2 U8883 ( .A1(a[16]), .A2(b[22]), .ZN(n7191) );
  INV_X4 U8884 ( .A(n7191), .ZN(n7189) );
  OAI21_X4 U8885 ( .B1(n7188), .B2(n7187), .A(n7186), .ZN(n7190) );
  NAND2_X2 U8886 ( .A1(n7189), .A2(n7190), .ZN(n7312) );
  INV_X4 U8887 ( .A(n7190), .ZN(n7192) );
  NAND2_X2 U8888 ( .A1(n7192), .A2(n7191), .ZN(n7311) );
  XNOR2_X2 U8889 ( .A(n7313), .B(n7193), .ZN(n7309) );
  NAND2_X2 U8890 ( .A1(a[17]), .A2(net246836), .ZN(n7201) );
  INV_X4 U8891 ( .A(n7201), .ZN(n7199) );
  INV_X4 U8892 ( .A(n7194), .ZN(n7195) );
  NAND2_X2 U8893 ( .A1(n7199), .A2(n7200), .ZN(n7308) );
  INV_X4 U8894 ( .A(n7200), .ZN(n7202) );
  NAND2_X2 U8895 ( .A1(n7202), .A2(n7201), .ZN(n7307) );
  NAND2_X2 U8896 ( .A1(n7308), .A2(n7307), .ZN(n7203) );
  XNOR2_X2 U8897 ( .A(n7309), .B(n7203), .ZN(n7304) );
  XNOR2_X2 U8898 ( .A(n7204), .B(n7304), .ZN(n7460) );
  XNOR2_X2 U8899 ( .A(n7460), .B(n7458), .ZN(n7211) );
  INV_X4 U8900 ( .A(n7205), .ZN(n7209) );
  INV_X4 U8901 ( .A(n7206), .ZN(n7207) );
  OAI21_X4 U8902 ( .B1(n7209), .B2(n7208), .A(n7207), .ZN(n7295) );
  NAND2_X2 U8903 ( .A1(n7209), .A2(n7208), .ZN(n7296) );
  NAND2_X2 U8904 ( .A1(n7295), .A2(n7296), .ZN(n7210) );
  XNOR2_X2 U8905 ( .A(n7211), .B(n7210), .ZN(n7290) );
  XNOR2_X2 U8906 ( .A(n7212), .B(n7290), .ZN(n7362) );
  XNOR2_X2 U8907 ( .A(n7213), .B(n7362), .ZN(n7375) );
  XNOR2_X2 U8908 ( .A(n7214), .B(n7375), .ZN(n7284) );
  INV_X4 U8909 ( .A(n7284), .ZN(n7215) );
  NAND2_X2 U8910 ( .A1(a[24]), .A2(b[14]), .ZN(n7274) );
  NAND2_X2 U8911 ( .A1(n7222), .A2(n7221), .ZN(n7276) );
  INV_X4 U8912 ( .A(net242906), .ZN(net242911) );
  NAND2_X2 U8913 ( .A1(b[13]), .A2(net246760), .ZN(net242908) );
  NAND2_X2 U8914 ( .A1(n7227), .A2(n7226), .ZN(net242910) );
  INV_X4 U8915 ( .A(net242910), .ZN(net242904) );
  INV_X4 U8916 ( .A(net242908), .ZN(net242907) );
  NAND2_X2 U8917 ( .A1(n7272), .A2(net242402), .ZN(n7228) );
  XNOR2_X2 U8918 ( .A(n4099), .B(n7228), .ZN(net242811) );
  INV_X4 U8919 ( .A(n7231), .ZN(n7230) );
  INV_X4 U8920 ( .A(net242879), .ZN(net242877) );
  NAND2_X2 U8921 ( .A1(b[8]), .A2(a[30]), .ZN(n7392) );
  XNOR2_X2 U8922 ( .A(n7393), .B(n7392), .ZN(n7234) );
  XNOR2_X2 U8923 ( .A(n7234), .B(n7396), .ZN(n7399) );
  NAND2_X2 U8924 ( .A1(net240782), .A2(a[7]), .ZN(n7235) );
  NAND2_X2 U8925 ( .A1(b[7]), .A2(n7236), .ZN(n7269) );
  NAND2_X2 U8926 ( .A1(net240913), .A2(net242655), .ZN(n7237) );
  NAND2_X2 U8927 ( .A1(n7237), .A2(n4550), .ZN(n7238) );
  NAND2_X2 U8928 ( .A1(n8784), .A2(n7239), .ZN(n7267) );
  NAND2_X2 U8929 ( .A1(n7242), .A2(n7240), .ZN(n7245) );
  INV_X4 U8930 ( .A(n7241), .ZN(n7244) );
  INV_X4 U8931 ( .A(n7242), .ZN(n7243) );
  AOI22_X2 U8932 ( .A1(n7245), .A2(n7244), .B1(n7243), .B2(a[8]), .ZN(n7410)
         );
  XNOR2_X2 U8933 ( .A(net246924), .B(b[7]), .ZN(n7408) );
  XNOR2_X2 U8934 ( .A(a[7]), .B(n7408), .ZN(n7246) );
  XNOR2_X2 U8935 ( .A(n7410), .B(n7246), .ZN(n7265) );
  NAND2_X2 U8936 ( .A1(n4558), .A2(n7658), .ZN(n7253) );
  NAND2_X2 U8937 ( .A1(n4562), .A2(n7247), .ZN(n7252) );
  NAND2_X2 U8938 ( .A1(n4554), .A2(n8118), .ZN(n7251) );
  AOI22_X2 U8939 ( .A1(net247082), .A2(a[23]), .B1(n8834), .B2(a[31]), .ZN(
        n7248) );
  OAI211_X2 U8940 ( .C1(net246958), .C2(n7409), .A(n7249), .B(n7248), .ZN(
        n8797) );
  NAND2_X2 U8941 ( .A1(n8797), .A2(n4565), .ZN(n7250) );
  NAND4_X2 U8942 ( .A1(n7253), .A2(n7252), .A3(n7251), .A4(n7250), .ZN(n7424)
         );
  NAND2_X2 U8943 ( .A1(n8318), .A2(n7424), .ZN(n7254) );
  AOI22_X2 U8944 ( .A1(n7256), .A2(n4564), .B1(n4557), .B2(n8111), .ZN(n7257)
         );
  OAI221_X2 U8945 ( .B1(n1323), .B2(n4533), .C1(n949), .C2(n8115), .A(n7257), 
        .ZN(n7258) );
  INV_X4 U8946 ( .A(n7258), .ZN(n7418) );
  NAND2_X2 U8947 ( .A1(net247002), .A2(a[7]), .ZN(n7262) );
  AOI21_X2 U8948 ( .B1(n4552), .B2(n7265), .A(n7264), .ZN(n7266) );
  NAND4_X2 U8949 ( .A1(n7269), .A2(n7268), .A3(n7267), .A4(n7266), .ZN(out[7])
         );
  NAND2_X2 U8950 ( .A1(net246772), .A2(b[10]), .ZN(n7440) );
  INV_X4 U8951 ( .A(n7440), .ZN(n7437) );
  NAND2_X2 U8952 ( .A1(b[11]), .A2(net246766), .ZN(n7442) );
  XNOR2_X2 U8953 ( .A(n7442), .B(n7438), .ZN(n7389) );
  NAND2_X2 U8954 ( .A1(net242821), .A2(net242819), .ZN(net242813) );
  NAND2_X2 U8955 ( .A1(b[12]), .A2(net246760), .ZN(n7450) );
  INV_X4 U8956 ( .A(net242819), .ZN(net242817) );
  NAND2_X2 U8957 ( .A1(n7450), .A2(net242812), .ZN(n7270) );
  NOR2_X4 U8958 ( .A1(n3909), .A2(n7270), .ZN(n7685) );
  INV_X4 U8959 ( .A(net242813), .ZN(net242581) );
  INV_X4 U8960 ( .A(net242812), .ZN(net242810) );
  NOR2_X4 U8961 ( .A1(n7271), .A2(n7685), .ZN(n7388) );
  XNOR2_X2 U8962 ( .A(n7273), .B(n3983), .ZN(n7386) );
  NAND2_X2 U8963 ( .A1(n7276), .A2(n7275), .ZN(n7277) );
  INV_X4 U8964 ( .A(n7277), .ZN(n7278) );
  NOR2_X4 U8965 ( .A1(n4091), .A2(n7278), .ZN(n7281) );
  OAI21_X4 U8966 ( .B1(n7281), .B2(n7280), .A(n7279), .ZN(n7611) );
  INV_X4 U8967 ( .A(n7611), .ZN(n7609) );
  NAND2_X2 U8968 ( .A1(a[23]), .A2(b[14]), .ZN(n7608) );
  INV_X4 U8969 ( .A(n7608), .ZN(n7612) );
  NAND2_X2 U8970 ( .A1(n7283), .A2(n7282), .ZN(n7285) );
  NAND2_X2 U8971 ( .A1(b[15]), .A2(a[22]), .ZN(n7605) );
  XNOR2_X2 U8972 ( .A(n7288), .B(n7605), .ZN(n7383) );
  NAND2_X2 U8973 ( .A1(n7290), .A2(n7289), .ZN(n7291) );
  OAI21_X4 U8974 ( .B1(n7293), .B2(n7292), .A(n7291), .ZN(n7574) );
  INV_X4 U8975 ( .A(n7574), .ZN(n7452) );
  NAND2_X2 U8976 ( .A1(a[19]), .A2(b[18]), .ZN(n7572) );
  NAND2_X2 U8977 ( .A1(b[17]), .A2(a[20]), .ZN(n7571) );
  XNOR2_X2 U8978 ( .A(n7572), .B(n7571), .ZN(n7294) );
  XNOR2_X2 U8979 ( .A(n7452), .B(n7294), .ZN(n7358) );
  INV_X4 U8980 ( .A(n7458), .ZN(n7299) );
  NAND2_X2 U8981 ( .A1(n7296), .A2(n7295), .ZN(n7297) );
  INV_X4 U8982 ( .A(n7297), .ZN(n7459) );
  NAND2_X2 U8983 ( .A1(n7299), .A2(n7298), .ZN(n7457) );
  NAND2_X2 U8984 ( .A1(a[17]), .A2(b[20]), .ZN(n7473) );
  INV_X4 U8985 ( .A(n7473), .ZN(n7306) );
  OAI21_X4 U8986 ( .B1(n7305), .B2(n4452), .A(n7303), .ZN(n7470) );
  XNOR2_X2 U8987 ( .A(n7306), .B(n7470), .ZN(n7356) );
  INV_X4 U8988 ( .A(n7307), .ZN(n7310) );
  NAND2_X2 U8989 ( .A1(n4578), .A2(net246836), .ZN(n7480) );
  NAND2_X2 U8990 ( .A1(a[15]), .A2(b[22]), .ZN(n7559) );
  INV_X4 U8991 ( .A(n7311), .ZN(n7314) );
  OAI21_X4 U8992 ( .B1(n7314), .B2(n7313), .A(n7312), .ZN(n7556) );
  XOR2_X2 U8993 ( .A(n7559), .B(n7556), .Z(n7355) );
  INV_X4 U8994 ( .A(n7315), .ZN(n7317) );
  NAND2_X2 U8995 ( .A1(n7317), .A2(n7316), .ZN(n7320) );
  NAND2_X2 U8996 ( .A1(a[7]), .A2(net248516), .ZN(n7484) );
  NAND3_X2 U8997 ( .A1(n7320), .A2(n7319), .A3(n3963), .ZN(n7485) );
  XNOR2_X2 U8998 ( .A(n7484), .B(n7721), .ZN(n7321) );
  XNOR2_X2 U8999 ( .A(n7485), .B(n7321), .ZN(n7490) );
  INV_X4 U9000 ( .A(n7322), .ZN(n7325) );
  OAI21_X4 U9001 ( .B1(n7325), .B2(n7324), .A(n7323), .ZN(n7491) );
  XOR2_X2 U9002 ( .A(n7490), .B(n7491), .Z(n7326) );
  NAND2_X2 U9003 ( .A1(a[8]), .A2(b[29]), .ZN(n7493) );
  XNOR2_X2 U9004 ( .A(n7326), .B(n7493), .ZN(n7501) );
  INV_X4 U9005 ( .A(n7327), .ZN(n7330) );
  OAI21_X4 U9006 ( .B1(n7330), .B2(n7329), .A(n7328), .ZN(n7500) );
  NAND2_X2 U9007 ( .A1(a[9]), .A2(net246880), .ZN(n7503) );
  INV_X4 U9008 ( .A(n7331), .ZN(n7334) );
  OAI21_X4 U9009 ( .B1(n7334), .B2(n7333), .A(n7332), .ZN(n7508) );
  NAND2_X2 U9010 ( .A1(a[10]), .A2(b[27]), .ZN(n7510) );
  INV_X4 U9011 ( .A(n7335), .ZN(n7338) );
  OAI21_X4 U9012 ( .B1(n7338), .B2(n7337), .A(n7336), .ZN(n7517) );
  XOR2_X2 U9013 ( .A(n7518), .B(n7517), .Z(n7339) );
  NAND2_X2 U9014 ( .A1(a[11]), .A2(b[26]), .ZN(n7520) );
  XNOR2_X2 U9015 ( .A(n7339), .B(n7520), .ZN(n7527) );
  INV_X4 U9016 ( .A(n7340), .ZN(n7343) );
  OAI21_X4 U9017 ( .B1(n7343), .B2(n7342), .A(n7341), .ZN(n7528) );
  NAND2_X2 U9018 ( .A1(a[12]), .A2(b[25]), .ZN(n7530) );
  INV_X4 U9019 ( .A(n7344), .ZN(n7347) );
  OAI21_X4 U9020 ( .B1(n7347), .B2(n7346), .A(n7345), .ZN(n7537) );
  XNOR2_X2 U9021 ( .A(n7538), .B(n7537), .ZN(n7349) );
  NAND2_X2 U9022 ( .A1(a[13]), .A2(b[24]), .ZN(n7540) );
  INV_X4 U9023 ( .A(n7540), .ZN(n7348) );
  XNOR2_X2 U9024 ( .A(n7349), .B(n7348), .ZN(n7548) );
  INV_X4 U9025 ( .A(n7350), .ZN(n7353) );
  OAI21_X4 U9026 ( .B1(n7353), .B2(n7352), .A(n7351), .ZN(n7547) );
  XNOR2_X2 U9027 ( .A(n7548), .B(n7547), .ZN(n7354) );
  XNOR2_X2 U9028 ( .A(n3976), .B(n7354), .ZN(n7557) );
  XNOR2_X2 U9029 ( .A(n7355), .B(n7557), .ZN(n7478) );
  XNOR2_X2 U9030 ( .A(n7356), .B(n7471), .ZN(n7463) );
  NAND2_X2 U9031 ( .A1(b[19]), .A2(a[18]), .ZN(n7466) );
  XNOR2_X2 U9032 ( .A(n7463), .B(n7466), .ZN(n7357) );
  XNOR2_X2 U9033 ( .A(n7464), .B(n7357), .ZN(n7573) );
  XNOR2_X2 U9034 ( .A(n7358), .B(n4468), .ZN(n7369) );
  NAND2_X2 U9035 ( .A1(n7359), .A2(n7082), .ZN(n7360) );
  AOI21_X4 U9036 ( .B1(n7367), .B2(n7366), .A(n7365), .ZN(n7368) );
  XNOR2_X2 U9037 ( .A(n7369), .B(n7368), .ZN(n7598) );
  NAND2_X2 U9038 ( .A1(a[21]), .A2(b[16]), .ZN(n7597) );
  XNOR2_X2 U9039 ( .A(n7370), .B(n7597), .ZN(n7381) );
  INV_X4 U9040 ( .A(n7373), .ZN(n7376) );
  NAND2_X2 U9041 ( .A1(n7376), .A2(n7374), .ZN(n7379) );
  INV_X4 U9042 ( .A(n7599), .ZN(n7380) );
  XNOR2_X2 U9043 ( .A(n7381), .B(n7380), .ZN(n7382) );
  XNOR2_X2 U9044 ( .A(n7383), .B(n7382), .ZN(n7610) );
  XNOR2_X2 U9045 ( .A(n7384), .B(n7610), .ZN(n7622) );
  XNOR2_X2 U9046 ( .A(n7386), .B(n7385), .ZN(n7684) );
  XNOR2_X2 U9047 ( .A(n7388), .B(n7387), .ZN(n7445) );
  XNOR2_X2 U9048 ( .A(n7391), .B(n7390), .ZN(net242611) );
  INV_X4 U9049 ( .A(n7392), .ZN(n7394) );
  OAI21_X4 U9050 ( .B1(n7396), .B2(n7397), .A(n7395), .ZN(net242379) );
  NAND2_X2 U9051 ( .A1(b[8]), .A2(net246786), .ZN(net242659) );
  INV_X4 U9052 ( .A(net242659), .ZN(net242378) );
  OAI22_X2 U9053 ( .A1(net242658), .A2(net242659), .B1(net242378), .B2(
        net242379), .ZN(n7398) );
  XNOR2_X2 U9054 ( .A(net248749), .B(n7398), .ZN(n7639) );
  INV_X4 U9055 ( .A(n7399), .ZN(n7400) );
  NAND2_X2 U9056 ( .A1(b[7]), .A2(a[30]), .ZN(n7635) );
  XNOR2_X2 U9057 ( .A(n7636), .B(n7635), .ZN(n7401) );
  XNOR2_X2 U9058 ( .A(n7639), .B(n7401), .ZN(n7436) );
  NAND2_X2 U9059 ( .A1(net240782), .A2(a[6]), .ZN(n7402) );
  NAND2_X2 U9060 ( .A1(b[6]), .A2(n7403), .ZN(n7435) );
  NAND2_X2 U9061 ( .A1(net240913), .A2(n7404), .ZN(n7405) );
  NAND2_X2 U9062 ( .A1(n7405), .A2(n4550), .ZN(n7406) );
  NAND2_X2 U9063 ( .A1(n8784), .A2(n7407), .ZN(n7433) );
  XNOR2_X2 U9064 ( .A(net246924), .B(b[6]), .ZN(n7649) );
  XNOR2_X2 U9065 ( .A(a[6]), .B(n7649), .ZN(n7414) );
  INV_X4 U9066 ( .A(n7408), .ZN(n7412) );
  NAND2_X2 U9067 ( .A1(n7410), .A2(n7409), .ZN(n7411) );
  OAI21_X4 U9068 ( .B1(n7413), .B2(n7412), .A(n7411), .ZN(n7650) );
  XNOR2_X2 U9069 ( .A(n7414), .B(n7650), .ZN(n7431) );
  NAND2_X2 U9070 ( .A1(n4562), .A2(n8845), .ZN(n7655) );
  AOI22_X2 U9071 ( .A1(n7415), .A2(n4564), .B1(n4557), .B2(n8314), .ZN(n7416)
         );
  OAI211_X2 U9072 ( .C1(n1386), .C2(n8115), .A(n7655), .B(n7416), .ZN(n7417)
         );
  INV_X4 U9073 ( .A(n7417), .ZN(n7668) );
  OAI22_X2 U9074 ( .A1(n7418), .A2(n4531), .B1(n7668), .B2(n4535), .ZN(n7427)
         );
  AOI22_X2 U9075 ( .A1(n4561), .A2(n7419), .B1(n4557), .B2(n7825), .ZN(n7423)
         );
  INV_X4 U9076 ( .A(n7424), .ZN(n7425) );
  OAI22_X2 U9077 ( .A1(n3986), .A2(n4537), .B1(n7425), .B2(n4539), .ZN(n7426)
         );
  NOR2_X2 U9078 ( .A1(n7427), .A2(n7426), .ZN(n7429) );
  NAND2_X2 U9079 ( .A1(net247002), .A2(a[6]), .ZN(n7428) );
  AOI21_X2 U9080 ( .B1(n4552), .B2(n7431), .A(n7430), .ZN(n7432) );
  NAND4_X2 U9081 ( .A1(n7435), .A2(n7434), .A3(n7433), .A4(n7432), .ZN(out[6])
         );
  NAND2_X2 U9082 ( .A1(b[6]), .A2(a[30]), .ZN(n7815) );
  XNOR2_X2 U9083 ( .A(n7816), .B(n7815), .ZN(n7642) );
  NAND2_X2 U9084 ( .A1(net246766), .A2(b[10]), .ZN(n7804) );
  XNOR2_X2 U9085 ( .A(n7438), .B(n7442), .ZN(n7439) );
  NAND2_X2 U9086 ( .A1(net242597), .A2(n7440), .ZN(n7799) );
  INV_X4 U9087 ( .A(n7442), .ZN(n7443) );
  INV_X4 U9088 ( .A(n7448), .ZN(n7446) );
  NAND2_X2 U9089 ( .A1(b[11]), .A2(net246760), .ZN(n7447) );
  INV_X4 U9090 ( .A(n7447), .ZN(n7449) );
  NAND2_X2 U9091 ( .A1(b[12]), .A2(net246754), .ZN(n7691) );
  XNOR2_X2 U9092 ( .A(n7451), .B(n7691), .ZN(n7633) );
  INV_X4 U9093 ( .A(n7572), .ZN(n7455) );
  INV_X4 U9094 ( .A(n7456), .ZN(n7768) );
  INV_X4 U9095 ( .A(n7457), .ZN(n7462) );
  NAND2_X2 U9096 ( .A1(n7464), .A2(n4462), .ZN(n7465) );
  OAI21_X4 U9097 ( .B1(n7467), .B2(n7466), .A(n7465), .ZN(n7712) );
  INV_X4 U9098 ( .A(n7712), .ZN(n7469) );
  NAND2_X2 U9099 ( .A1(a[17]), .A2(b[19]), .ZN(n7468) );
  INV_X4 U9100 ( .A(n7468), .ZN(n7713) );
  AOI22_X2 U9101 ( .A1(n7469), .A2(n7468), .B1(n7713), .B2(n7712), .ZN(n7569)
         );
  AOI21_X4 U9102 ( .B1(a[16]), .B2(b[20]), .A(n7475), .ZN(n7717) );
  NAND2_X2 U9103 ( .A1(n4578), .A2(n7475), .ZN(n7716) );
  INV_X4 U9104 ( .A(n7716), .ZN(n7476) );
  NOR2_X4 U9105 ( .A1(n7717), .A2(n7476), .ZN(n7567) );
  OAI21_X4 U9106 ( .B1(n7481), .B2(n7480), .A(n7479), .ZN(n7482) );
  AOI21_X4 U9107 ( .B1(a[15]), .B2(net246836), .A(n7482), .ZN(n7764) );
  NAND2_X2 U9108 ( .A1(a[15]), .A2(n7482), .ZN(n7762) );
  INV_X4 U9109 ( .A(n7762), .ZN(n7483) );
  NOR2_X4 U9110 ( .A1(n7764), .A2(n7483), .ZN(n7566) );
  INV_X4 U9111 ( .A(n7484), .ZN(n7486) );
  NAND2_X2 U9112 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  OAI21_X4 U9113 ( .B1(n7488), .B2(n7721), .A(n7487), .ZN(n7718) );
  XOR2_X2 U9114 ( .A(n7719), .B(n7718), .Z(n7489) );
  NAND2_X2 U9115 ( .A1(a[6]), .A2(net248517), .ZN(n7720) );
  XNOR2_X2 U9116 ( .A(n7489), .B(n7720), .ZN(n7726) );
  NAND2_X2 U9117 ( .A1(a[7]), .A2(b[29]), .ZN(n7497) );
  INV_X4 U9118 ( .A(n7497), .ZN(n7495) );
  NAND2_X2 U9119 ( .A1(n7491), .A2(n7490), .ZN(n7492) );
  OAI21_X4 U9120 ( .B1(n7494), .B2(n7493), .A(n7492), .ZN(n7496) );
  NAND2_X2 U9121 ( .A1(n7495), .A2(n7496), .ZN(n7725) );
  INV_X4 U9122 ( .A(n7496), .ZN(n7498) );
  NAND2_X2 U9123 ( .A1(n7498), .A2(n7497), .ZN(n7724) );
  NAND2_X2 U9124 ( .A1(n7725), .A2(n7724), .ZN(n7499) );
  XNOR2_X2 U9125 ( .A(n7726), .B(n7499), .ZN(n7730) );
  NAND2_X2 U9126 ( .A1(n3970), .A2(n7505), .ZN(n7729) );
  NAND2_X2 U9127 ( .A1(n7729), .A2(n7728), .ZN(n7506) );
  XNOR2_X2 U9128 ( .A(n7730), .B(n7506), .ZN(n7734) );
  NAND2_X2 U9129 ( .A1(a[9]), .A2(b[27]), .ZN(n7514) );
  INV_X4 U9130 ( .A(n7514), .ZN(n7512) );
  NAND2_X2 U9131 ( .A1(n7508), .A2(n7507), .ZN(n7509) );
  OAI21_X4 U9132 ( .B1(n7511), .B2(n7510), .A(n7509), .ZN(n7513) );
  NAND2_X2 U9133 ( .A1(n7512), .A2(n7513), .ZN(n7733) );
  INV_X4 U9134 ( .A(n7513), .ZN(n7515) );
  NAND2_X2 U9135 ( .A1(n7515), .A2(n7514), .ZN(n7732) );
  NAND2_X2 U9136 ( .A1(n7733), .A2(n7732), .ZN(n7516) );
  XNOR2_X2 U9137 ( .A(n7734), .B(n7516), .ZN(n7739) );
  NAND2_X2 U9138 ( .A1(a[10]), .A2(b[26]), .ZN(n7524) );
  INV_X4 U9139 ( .A(n7524), .ZN(n7522) );
  NAND2_X2 U9140 ( .A1(n4433), .A2(n7517), .ZN(n7519) );
  OAI21_X4 U9141 ( .B1(n7521), .B2(n7520), .A(n7519), .ZN(n7523) );
  NAND2_X2 U9142 ( .A1(n7522), .A2(n7523), .ZN(n7738) );
  INV_X4 U9143 ( .A(n7523), .ZN(n7525) );
  NAND2_X2 U9144 ( .A1(n7525), .A2(n7524), .ZN(n7737) );
  NAND2_X2 U9145 ( .A1(n7738), .A2(n7737), .ZN(n7526) );
  XNOR2_X2 U9146 ( .A(n7739), .B(n7526), .ZN(n7744) );
  NAND2_X2 U9147 ( .A1(a[11]), .A2(b[25]), .ZN(n7534) );
  INV_X4 U9148 ( .A(n7534), .ZN(n7532) );
  NAND2_X2 U9149 ( .A1(n7528), .A2(n7527), .ZN(n7529) );
  OAI21_X4 U9150 ( .B1(n7531), .B2(n7530), .A(n7529), .ZN(n7533) );
  NAND2_X2 U9151 ( .A1(n7532), .A2(n7533), .ZN(n7743) );
  INV_X4 U9152 ( .A(n7533), .ZN(n7535) );
  NAND2_X2 U9153 ( .A1(n7535), .A2(n7534), .ZN(n7742) );
  NAND2_X2 U9154 ( .A1(n7743), .A2(n7742), .ZN(n7536) );
  XNOR2_X2 U9155 ( .A(n7744), .B(n7536), .ZN(n7748) );
  NAND2_X2 U9156 ( .A1(a[12]), .A2(b[24]), .ZN(n7544) );
  INV_X4 U9157 ( .A(n7544), .ZN(n7542) );
  NAND2_X2 U9158 ( .A1(n7538), .A2(n7537), .ZN(n7539) );
  OAI21_X4 U9159 ( .B1(n7541), .B2(n7540), .A(n7539), .ZN(n7543) );
  NAND2_X2 U9160 ( .A1(n7542), .A2(n7543), .ZN(n7747) );
  INV_X4 U9161 ( .A(n7543), .ZN(n7545) );
  NAND2_X2 U9162 ( .A1(n7545), .A2(n7544), .ZN(n7746) );
  NAND2_X2 U9163 ( .A1(n7747), .A2(n7746), .ZN(n7546) );
  XNOR2_X2 U9164 ( .A(n7748), .B(n7546), .ZN(n7753) );
  NAND2_X2 U9165 ( .A1(a[13]), .A2(b[23]), .ZN(n7553) );
  INV_X4 U9166 ( .A(n7553), .ZN(n7551) );
  NAND2_X2 U9167 ( .A1(n7547), .A2(n7548), .ZN(n7550) );
  NAND2_X2 U9168 ( .A1(n7550), .A2(n7549), .ZN(n7552) );
  NAND2_X2 U9169 ( .A1(n7551), .A2(n7552), .ZN(n7752) );
  INV_X4 U9170 ( .A(n7552), .ZN(n7554) );
  NAND2_X2 U9171 ( .A1(n7554), .A2(n7553), .ZN(n7751) );
  NAND2_X2 U9172 ( .A1(n7752), .A2(n7751), .ZN(n7555) );
  XNOR2_X2 U9173 ( .A(n7753), .B(n7555), .ZN(n7758) );
  NAND2_X2 U9174 ( .A1(a[14]), .A2(b[22]), .ZN(n7563) );
  INV_X4 U9175 ( .A(n7563), .ZN(n7561) );
  OAI21_X4 U9176 ( .B1(n7560), .B2(n7559), .A(n7558), .ZN(n7562) );
  NAND2_X2 U9177 ( .A1(n7561), .A2(n7562), .ZN(n7757) );
  INV_X4 U9178 ( .A(n7562), .ZN(n7564) );
  NAND2_X2 U9179 ( .A1(n7564), .A2(n7563), .ZN(n7756) );
  NAND2_X2 U9180 ( .A1(n7757), .A2(n7756), .ZN(n7565) );
  XNOR2_X2 U9181 ( .A(n7758), .B(n7565), .ZN(n7763) );
  INV_X4 U9182 ( .A(n7711), .ZN(n7568) );
  XNOR2_X2 U9183 ( .A(n7569), .B(n7568), .ZN(n7769) );
  XNOR2_X2 U9184 ( .A(n7769), .B(n7767), .ZN(n7570) );
  XNOR2_X2 U9185 ( .A(n7768), .B(n7570), .ZN(n7774) );
  NAND2_X2 U9186 ( .A1(b[17]), .A2(a[19]), .ZN(n7584) );
  INV_X4 U9187 ( .A(n7584), .ZN(n7582) );
  INV_X4 U9188 ( .A(n7571), .ZN(n7576) );
  NAND2_X2 U9189 ( .A1(n7576), .A2(n7577), .ZN(n7581) );
  XNOR2_X2 U9190 ( .A(n7573), .B(n7572), .ZN(n7575) );
  XNOR2_X2 U9191 ( .A(n7575), .B(n7574), .ZN(n7578) );
  NAND2_X2 U9192 ( .A1(n7576), .A2(n7578), .ZN(n7580) );
  NAND2_X2 U9193 ( .A1(n7578), .A2(n7577), .ZN(n7579) );
  NAND3_X4 U9194 ( .A1(n7581), .A2(n7580), .A3(n7579), .ZN(n7583) );
  NAND2_X2 U9195 ( .A1(n7582), .A2(n7583), .ZN(n7773) );
  INV_X4 U9196 ( .A(n7583), .ZN(n7585) );
  NAND2_X2 U9197 ( .A1(n7585), .A2(n7584), .ZN(n7772) );
  NAND2_X2 U9198 ( .A1(n7773), .A2(n7772), .ZN(n7586) );
  XNOR2_X2 U9199 ( .A(n7774), .B(n7586), .ZN(n7708) );
  NAND2_X2 U9200 ( .A1(n7588), .A2(n7587), .ZN(n7591) );
  INV_X4 U9201 ( .A(n7591), .ZN(n7590) );
  NAND2_X2 U9202 ( .A1(a[20]), .A2(b[16]), .ZN(n7592) );
  INV_X4 U9203 ( .A(n7592), .ZN(n7589) );
  NAND2_X2 U9204 ( .A1(n7590), .A2(n7589), .ZN(n7707) );
  NAND2_X2 U9205 ( .A1(n7592), .A2(n7591), .ZN(n7706) );
  XNOR2_X2 U9206 ( .A(n7594), .B(n7593), .ZN(n7785) );
  INV_X4 U9207 ( .A(n7288), .ZN(n7601) );
  XNOR2_X2 U9208 ( .A(n7600), .B(n7599), .ZN(n7602) );
  NAND2_X2 U9209 ( .A1(n7601), .A2(n7602), .ZN(n7781) );
  INV_X4 U9210 ( .A(n7781), .ZN(n7606) );
  INV_X4 U9211 ( .A(n7605), .ZN(n7782) );
  NAND2_X2 U9212 ( .A1(n7782), .A2(a[21]), .ZN(n7604) );
  NAND2_X2 U9213 ( .A1(b[15]), .A2(a[21]), .ZN(n7779) );
  INV_X4 U9214 ( .A(n7602), .ZN(n7603) );
  OAI211_X2 U9215 ( .C1(n7606), .C2(n7605), .A(n7779), .B(n7780), .ZN(n7697)
         );
  XNOR2_X2 U9216 ( .A(n4463), .B(n7607), .ZN(n7619) );
  NAND2_X2 U9217 ( .A1(a[22]), .A2(b[14]), .ZN(n7703) );
  INV_X4 U9218 ( .A(n7703), .ZN(n7615) );
  NAND3_X4 U9219 ( .A1(n7617), .A2(n7616), .A3(n7615), .ZN(n8054) );
  INV_X4 U9220 ( .A(n7616), .ZN(n7704) );
  OAI21_X4 U9221 ( .B1(n7704), .B2(n4040), .A(n7703), .ZN(n7618) );
  NAND2_X2 U9222 ( .A1(n8054), .A2(n7618), .ZN(n7699) );
  XNOR2_X2 U9223 ( .A(n7619), .B(n7699), .ZN(n7687) );
  INV_X4 U9224 ( .A(n7687), .ZN(n7631) );
  NAND2_X2 U9225 ( .A1(n3983), .A2(n7621), .ZN(n7624) );
  NAND2_X2 U9226 ( .A1(n7622), .A2(n7621), .ZN(n7623) );
  NAND3_X2 U9227 ( .A1(n7625), .A2(n7624), .A3(n7623), .ZN(n7628) );
  INV_X4 U9228 ( .A(n7628), .ZN(n7626) );
  NAND2_X2 U9229 ( .A1(b[13]), .A2(a[23]), .ZN(n7627) );
  INV_X4 U9230 ( .A(n7627), .ZN(n7629) );
  NAND2_X2 U9231 ( .A1(n7629), .A2(n7628), .ZN(n8068) );
  NAND2_X2 U9232 ( .A1(n7700), .A2(n8068), .ZN(n7630) );
  XNOR2_X2 U9233 ( .A(n7631), .B(n7630), .ZN(n7632) );
  XNOR2_X2 U9234 ( .A(n7634), .B(n7796), .ZN(net242385) );
  NAND2_X2 U9235 ( .A1(net242378), .A2(net242379), .ZN(net242316) );
  INV_X4 U9236 ( .A(net242316), .ZN(net242311) );
  INV_X4 U9237 ( .A(n7635), .ZN(n7637) );
  OAI21_X4 U9238 ( .B1(n7639), .B2(n7640), .A(n7638), .ZN(net242324) );
  NAND2_X2 U9239 ( .A1(b[7]), .A2(net246788), .ZN(net242367) );
  XNOR2_X2 U9240 ( .A(net248078), .B(net242366), .ZN(n7862) );
  XNOR2_X2 U9241 ( .A(n7641), .B(n7642), .ZN(n7820) );
  NAND2_X2 U9242 ( .A1(net240782), .A2(a[5]), .ZN(n7643) );
  NAND2_X2 U9243 ( .A1(n7644), .A2(b[5]), .ZN(n7678) );
  NAND2_X2 U9244 ( .A1(net240913), .A2(net242361), .ZN(n7645) );
  NAND2_X2 U9245 ( .A1(n7645), .A2(n4550), .ZN(n7646) );
  NAND2_X2 U9246 ( .A1(n8784), .A2(n7647), .ZN(n7676) );
  NAND2_X2 U9247 ( .A1(n7650), .A2(n7648), .ZN(n7653) );
  INV_X4 U9248 ( .A(n7649), .ZN(n7652) );
  INV_X4 U9249 ( .A(n7650), .ZN(n7651) );
  AOI22_X2 U9250 ( .A1(n7653), .A2(n7652), .B1(n7651), .B2(a[6]), .ZN(n7843)
         );
  XNOR2_X2 U9251 ( .A(net246924), .B(b[5]), .ZN(n7841) );
  XNOR2_X2 U9252 ( .A(a[5]), .B(n7841), .ZN(n7654) );
  XNOR2_X2 U9253 ( .A(n7843), .B(n7654), .ZN(n7674) );
  INV_X4 U9254 ( .A(n7655), .ZN(n7656) );
  OAI221_X2 U9255 ( .B1(n1323), .B2(n8832), .C1(n949), .C2(n4566), .A(n7657), 
        .ZN(n7836) );
  INV_X4 U9256 ( .A(n7836), .ZN(n7667) );
  NAND2_X2 U9257 ( .A1(n4555), .A2(n8797), .ZN(n7665) );
  NAND2_X2 U9258 ( .A1(n4562), .A2(n7658), .ZN(n7664) );
  NAND2_X2 U9259 ( .A1(n4559), .A2(n8118), .ZN(n7663) );
  NAND2_X2 U9260 ( .A1(net246962), .A2(a[5]), .ZN(n7661) );
  AOI22_X2 U9261 ( .A1(net247082), .A2(a[21]), .B1(n8834), .B2(net246788), 
        .ZN(n7659) );
  NAND3_X2 U9262 ( .A1(n7661), .A2(n7660), .A3(n7659), .ZN(n8795) );
  NAND2_X2 U9263 ( .A1(n8795), .A2(n4565), .ZN(n7662) );
  NAND4_X2 U9264 ( .A1(n7665), .A2(n7664), .A3(n7663), .A4(n7662), .ZN(n7833)
         );
  NAND2_X2 U9265 ( .A1(n8318), .A2(n7833), .ZN(n7666) );
  OAI22_X2 U9266 ( .A1(n7668), .A2(n4531), .B1(n3986), .B2(n4539), .ZN(n7669)
         );
  NAND2_X2 U9267 ( .A1(net247002), .A2(a[5]), .ZN(n7671) );
  AOI21_X2 U9268 ( .B1(n4552), .B2(n7674), .A(n7673), .ZN(n7675) );
  NAND4_X2 U9269 ( .A1(n7678), .A2(n7677), .A3(n7676), .A4(n7675), .ZN(out[5])
         );
  NAND2_X2 U9270 ( .A1(b[6]), .A2(net246788), .ZN(n7869) );
  XNOR2_X2 U9271 ( .A(n7869), .B(net241613), .ZN(net242322) );
  NAND2_X2 U9272 ( .A1(net246772), .A2(b[8]), .ZN(n7681) );
  INV_X4 U9273 ( .A(n7681), .ZN(n7877) );
  OAI21_X4 U9274 ( .B1(n7680), .B2(net242309), .A(net242310), .ZN(n7876) );
  XNOR2_X2 U9275 ( .A(n7683), .B(net241760), .ZN(net242153) );
  NAND2_X2 U9276 ( .A1(b[12]), .A2(a[23]), .ZN(n7882) );
  NAND2_X2 U9277 ( .A1(n7686), .A2(n7691), .ZN(n7690) );
  NAND2_X2 U9278 ( .A1(n8068), .A2(n7700), .ZN(n7688) );
  XNOR2_X2 U9279 ( .A(n7688), .B(n7687), .ZN(n7689) );
  INV_X4 U9280 ( .A(n7691), .ZN(n7693) );
  XNOR2_X2 U9281 ( .A(n7882), .B(n7694), .ZN(n7794) );
  INV_X4 U9282 ( .A(n7695), .ZN(n7696) );
  XNOR2_X2 U9283 ( .A(n7698), .B(n7785), .ZN(n8053) );
  XNOR2_X2 U9284 ( .A(n4400), .B(n7699), .ZN(n7701) );
  NAND2_X2 U9285 ( .A1(n7701), .A2(n7700), .ZN(n8069) );
  NAND2_X2 U9286 ( .A1(b[13]), .A2(a[22]), .ZN(n8067) );
  XNOR2_X2 U9287 ( .A(n7702), .B(n8067), .ZN(n7793) );
  INV_X4 U9288 ( .A(n8054), .ZN(n7705) );
  INV_X4 U9289 ( .A(n7706), .ZN(n7709) );
  OAI21_X4 U9290 ( .B1(n7709), .B2(n7708), .A(n7707), .ZN(n8033) );
  NAND2_X2 U9291 ( .A1(a[19]), .A2(b[16]), .ZN(n8032) );
  NAND2_X2 U9292 ( .A1(b[15]), .A2(a[20]), .ZN(n8031) );
  XNOR2_X2 U9293 ( .A(n8032), .B(n8031), .ZN(n7710) );
  XNOR2_X2 U9294 ( .A(n8033), .B(n7710), .ZN(n7777) );
  OAI21_X4 U9295 ( .B1(n7713), .B2(n7712), .A(n7711), .ZN(n7715) );
  NAND2_X2 U9296 ( .A1(n7713), .A2(n7712), .ZN(n7714) );
  NAND2_X2 U9297 ( .A1(n7715), .A2(n7714), .ZN(n7895) );
  NAND2_X2 U9298 ( .A1(a[15]), .A2(b[20]), .ZN(n7905) );
  OAI21_X4 U9299 ( .B1(n7717), .B2(n3946), .A(n7716), .ZN(n7902) );
  XOR2_X2 U9300 ( .A(n7905), .B(n7902), .Z(n7765) );
  INV_X4 U9301 ( .A(n7718), .ZN(n7722) );
  NAND2_X2 U9302 ( .A1(a[5]), .A2(net246902), .ZN(n7909) );
  OAI21_X4 U9303 ( .B1(n7722), .B2(n3940), .A(n3973), .ZN(n7910) );
  XNOR2_X2 U9304 ( .A(n7909), .B(n8197), .ZN(n7723) );
  XNOR2_X2 U9305 ( .A(n7910), .B(n7723), .ZN(n7916) );
  INV_X4 U9306 ( .A(n7724), .ZN(n7727) );
  OAI21_X4 U9307 ( .B1(n7727), .B2(n7726), .A(n7725), .ZN(n7917) );
  NAND2_X2 U9308 ( .A1(a[6]), .A2(b[29]), .ZN(n7919) );
  OAI21_X4 U9309 ( .B1(n4445), .B2(n7730), .A(n7729), .ZN(n7926) );
  XOR2_X2 U9310 ( .A(n7927), .B(n7926), .Z(n7731) );
  NAND2_X2 U9311 ( .A1(a[7]), .A2(net246880), .ZN(n7929) );
  XNOR2_X2 U9312 ( .A(n7731), .B(n7929), .ZN(n7936) );
  INV_X4 U9313 ( .A(n7732), .ZN(n7735) );
  OAI21_X4 U9314 ( .B1(n7735), .B2(n7734), .A(n7733), .ZN(n7937) );
  XOR2_X2 U9315 ( .A(n7936), .B(n7937), .Z(n7736) );
  NAND2_X2 U9316 ( .A1(a[8]), .A2(b[27]), .ZN(n7939) );
  XNOR2_X2 U9317 ( .A(n7736), .B(n7939), .ZN(n7947) );
  INV_X4 U9318 ( .A(n7737), .ZN(n7740) );
  OAI21_X4 U9319 ( .B1(n7740), .B2(n7739), .A(n7738), .ZN(n7946) );
  XOR2_X2 U9320 ( .A(n7947), .B(n7946), .Z(n7741) );
  NAND2_X2 U9321 ( .A1(a[9]), .A2(b[26]), .ZN(n7949) );
  XNOR2_X2 U9322 ( .A(n7741), .B(n7949), .ZN(n7956) );
  INV_X4 U9323 ( .A(n7742), .ZN(n7745) );
  OAI21_X4 U9324 ( .B1(n7745), .B2(n7744), .A(n7743), .ZN(n7957) );
  NAND2_X2 U9325 ( .A1(a[10]), .A2(b[25]), .ZN(n7959) );
  INV_X4 U9326 ( .A(n7746), .ZN(n7749) );
  OAI21_X4 U9327 ( .B1(n7749), .B2(n7748), .A(n7747), .ZN(n7966) );
  XOR2_X2 U9328 ( .A(n7967), .B(n7966), .Z(n7750) );
  NAND2_X2 U9329 ( .A1(a[11]), .A2(b[24]), .ZN(n7969) );
  XNOR2_X2 U9330 ( .A(n7750), .B(n7969), .ZN(n7976) );
  INV_X4 U9331 ( .A(n7751), .ZN(n7754) );
  OAI21_X4 U9332 ( .B1(n7754), .B2(n7753), .A(n7752), .ZN(n7977) );
  XOR2_X2 U9333 ( .A(n7976), .B(n7977), .Z(n7755) );
  NAND2_X2 U9334 ( .A1(a[12]), .A2(b[23]), .ZN(n7979) );
  XNOR2_X2 U9335 ( .A(n7755), .B(n7979), .ZN(n7987) );
  INV_X4 U9336 ( .A(n7756), .ZN(n7759) );
  OAI21_X4 U9337 ( .B1(n7759), .B2(n7758), .A(n7757), .ZN(n7986) );
  XNOR2_X2 U9338 ( .A(n7987), .B(n7986), .ZN(n7761) );
  NAND2_X2 U9339 ( .A1(a[13]), .A2(b[22]), .ZN(n7989) );
  INV_X4 U9340 ( .A(n7989), .ZN(n7760) );
  XNOR2_X2 U9341 ( .A(n7761), .B(n7760), .ZN(n7996) );
  NAND2_X2 U9342 ( .A1(a[14]), .A2(net246836), .ZN(n7999) );
  OAI21_X4 U9343 ( .B1(n7764), .B2(n7763), .A(n7762), .ZN(n7997) );
  XNOR2_X2 U9344 ( .A(n7765), .B(n7903), .ZN(n7894) );
  NAND2_X2 U9345 ( .A1(n4578), .A2(b[19]), .ZN(n7893) );
  XNOR2_X2 U9346 ( .A(n7894), .B(n7893), .ZN(n7766) );
  XNOR2_X2 U9347 ( .A(n7895), .B(n7766), .ZN(n8009) );
  NAND2_X2 U9348 ( .A1(a[17]), .A2(b[18]), .ZN(n8010) );
  INV_X4 U9349 ( .A(n7767), .ZN(n7770) );
  OAI21_X4 U9350 ( .B1(n7770), .B2(n4444), .A(n7768), .ZN(n8011) );
  NAND2_X2 U9351 ( .A1(n7770), .A2(n4444), .ZN(n8012) );
  OAI21_X4 U9352 ( .B1(n7775), .B2(n7774), .A(n7773), .ZN(n8024) );
  NAND2_X2 U9353 ( .A1(b[17]), .A2(a[18]), .ZN(n8022) );
  XNOR2_X2 U9354 ( .A(n8024), .B(n8022), .ZN(n7776) );
  XNOR2_X2 U9355 ( .A(n8025), .B(n7776), .ZN(n8034) );
  XNOR2_X2 U9356 ( .A(n8034), .B(n7777), .ZN(n8048) );
  XNOR2_X2 U9357 ( .A(n7778), .B(n8048), .ZN(n7792) );
  INV_X4 U9358 ( .A(n7779), .ZN(n7784) );
  INV_X4 U9359 ( .A(n7780), .ZN(n7787) );
  NAND2_X2 U9360 ( .A1(n7782), .A2(n7781), .ZN(n7783) );
  INV_X4 U9361 ( .A(n7783), .ZN(n7786) );
  NOR3_X4 U9362 ( .A1(n7784), .A2(n7787), .A3(n7786), .ZN(n7790) );
  INV_X4 U9363 ( .A(n4463), .ZN(n7789) );
  OAI21_X4 U9364 ( .B1(n7787), .B2(n7786), .A(a[21]), .ZN(n7788) );
  OAI21_X4 U9365 ( .B1(n7790), .B2(n7789), .A(n7788), .ZN(n8037) );
  INV_X4 U9366 ( .A(n8037), .ZN(n8049) );
  NAND2_X2 U9367 ( .A1(a[21]), .A2(b[14]), .ZN(n8060) );
  XNOR2_X2 U9368 ( .A(n8049), .B(n8060), .ZN(n7791) );
  XNOR2_X2 U9369 ( .A(n7792), .B(n7791), .ZN(n8071) );
  XNOR2_X2 U9370 ( .A(n7793), .B(n8071), .ZN(n7878) );
  XNOR2_X2 U9371 ( .A(n7794), .B(n7878), .ZN(n8080) );
  NAND2_X2 U9372 ( .A1(b[11]), .A2(net246754), .ZN(n8084) );
  INV_X4 U9373 ( .A(n8084), .ZN(n8086) );
  XNOR2_X2 U9374 ( .A(n7797), .B(n8086), .ZN(n7798) );
  XNOR2_X2 U9375 ( .A(n7798), .B(n8080), .ZN(n8096) );
  NAND2_X2 U9376 ( .A1(n7799), .A2(n7800), .ZN(n7803) );
  INV_X4 U9377 ( .A(n7811), .ZN(n7810) );
  INV_X4 U9378 ( .A(n7813), .ZN(n7809) );
  INV_X4 U9379 ( .A(n7803), .ZN(n7806) );
  INV_X4 U9380 ( .A(n7804), .ZN(n7805) );
  INV_X4 U9381 ( .A(n7807), .ZN(n7812) );
  NOR2_X4 U9382 ( .A1(n7812), .A2(n3980), .ZN(n7808) );
  OAI21_X4 U9383 ( .B1(n7810), .B2(n7809), .A(n7808), .ZN(n8095) );
  XNOR2_X2 U9384 ( .A(n8096), .B(n7814), .ZN(net241826) );
  XNOR2_X2 U9385 ( .A(net242151), .B(net242097), .ZN(n7819) );
  INV_X4 U9386 ( .A(n7863), .ZN(n7866) );
  INV_X4 U9387 ( .A(n7815), .ZN(n7818) );
  NAND2_X2 U9388 ( .A1(n7818), .A2(n7817), .ZN(n7861) );
  XNOR2_X2 U9389 ( .A(n7819), .B(n7868), .ZN(n7855) );
  NAND2_X2 U9390 ( .A1(b[5]), .A2(a[30]), .ZN(n7856) );
  XNOR2_X2 U9391 ( .A(n7855), .B(n7821), .ZN(n7823) );
  NAND2_X2 U9392 ( .A1(net240913), .A2(net242110), .ZN(n7824) );
  NAND2_X2 U9393 ( .A1(n7824), .A2(n4550), .ZN(n7840) );
  INV_X4 U9394 ( .A(n7825), .ZN(n7831) );
  INV_X4 U9395 ( .A(n8303), .ZN(n7829) );
  AOI22_X2 U9396 ( .A1(net247082), .A2(a[20]), .B1(n8834), .B2(a[28]), .ZN(
        n7826) );
  OAI211_X2 U9397 ( .C1(net246958), .C2(n8130), .A(n7827), .B(n7826), .ZN(
        n8831) );
  AOI22_X2 U9398 ( .A1(n8831), .A2(n4564), .B1(n4557), .B2(n8305), .ZN(n7828)
         );
  OAI221_X2 U9399 ( .B1(n7831), .B2(n4533), .C1(n7829), .C2(n8115), .A(n7828), 
        .ZN(n8110) );
  AOI22_X2 U9400 ( .A1(n8318), .A2(n8110), .B1(n8125), .B2(n8109), .ZN(n7838)
         );
  INV_X4 U9401 ( .A(n7833), .ZN(n7834) );
  AOI21_X2 U9402 ( .B1(n8842), .B2(n7836), .A(n7835), .ZN(n7837) );
  XNOR2_X2 U9403 ( .A(net246924), .B(b[4]), .ZN(n8131) );
  XNOR2_X2 U9404 ( .A(a[4]), .B(n8131), .ZN(n7847) );
  INV_X4 U9405 ( .A(n7841), .ZN(n7845) );
  NAND2_X2 U9406 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  OAI21_X4 U9407 ( .B1(n7846), .B2(n7845), .A(n7844), .ZN(n8132) );
  XNOR2_X2 U9408 ( .A(n7847), .B(n8132), .ZN(n7851) );
  NAND2_X2 U9409 ( .A1(n8784), .A2(n7848), .ZN(n7849) );
  AOI21_X2 U9410 ( .B1(n4552), .B2(n7851), .A(n7850), .ZN(n7852) );
  OAI211_X2 U9411 ( .C1(n7854), .C2(net242110), .A(n7852), .B(n7853), .ZN(
        out[4]) );
  NAND2_X2 U9412 ( .A1(b[5]), .A2(net246786), .ZN(net241579) );
  NAND2_X2 U9413 ( .A1(n7856), .A2(n7857), .ZN(n7858) );
  NAND2_X2 U9414 ( .A1(n7858), .A2(n8273), .ZN(net242103) );
  INV_X4 U9415 ( .A(n7858), .ZN(n8274) );
  INV_X4 U9416 ( .A(net242102), .ZN(net242099) );
  XNOR2_X2 U9417 ( .A(n7860), .B(net242097), .ZN(net242095) );
  INV_X4 U9418 ( .A(net242095), .ZN(net242079) );
  INV_X4 U9419 ( .A(n7869), .ZN(n7864) );
  OAI21_X4 U9420 ( .B1(n7866), .B2(n3910), .A(n7869), .ZN(n7871) );
  OAI21_X4 U9421 ( .B1(net242079), .B2(n7867), .A(n7871), .ZN(net241770) );
  NAND2_X2 U9422 ( .A1(b[6]), .A2(a[28]), .ZN(net241771) );
  INV_X4 U9423 ( .A(n7868), .ZN(n7870) );
  INV_X4 U9424 ( .A(n7871), .ZN(n7872) );
  NOR2_X4 U9425 ( .A1(n7872), .A2(net241771), .ZN(net242080) );
  NAND2_X2 U9426 ( .A1(net246766), .A2(b[8]), .ZN(n8269) );
  NOR2_X4 U9427 ( .A1(net242066), .A2(net242067), .ZN(n7873) );
  XNOR2_X2 U9428 ( .A(n7873), .B(net241760), .ZN(n7874) );
  XNOR2_X2 U9429 ( .A(n7874), .B(net241826), .ZN(n7875) );
  NAND2_X2 U9430 ( .A1(b[12]), .A2(a[22]), .ZN(n7890) );
  INV_X4 U9431 ( .A(n7890), .ZN(n7888) );
  INV_X4 U9432 ( .A(n7882), .ZN(n7879) );
  INV_X4 U9433 ( .A(n7878), .ZN(n7884) );
  NAND2_X2 U9434 ( .A1(n7879), .A2(n7884), .ZN(n7887) );
  NAND2_X2 U9435 ( .A1(n7883), .A2(n7879), .ZN(n7886) );
  NAND2_X2 U9436 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  NAND2_X2 U9437 ( .A1(n4425), .A2(n7888), .ZN(n8157) );
  INV_X4 U9438 ( .A(n7889), .ZN(n7891) );
  NAND2_X2 U9439 ( .A1(n7891), .A2(n7890), .ZN(n8156) );
  NAND2_X2 U9440 ( .A1(n8157), .A2(n8156), .ZN(n7892) );
  INV_X4 U9441 ( .A(n7893), .ZN(n7896) );
  NAND2_X2 U9442 ( .A1(n7896), .A2(n7895), .ZN(n7897) );
  NAND3_X2 U9443 ( .A1(n7899), .A2(n7898), .A3(n7897), .ZN(n7900) );
  AOI21_X4 U9444 ( .B1(a[15]), .B2(b[19]), .A(n7900), .ZN(n8193) );
  NAND2_X2 U9445 ( .A1(a[15]), .A2(n7900), .ZN(n8191) );
  INV_X4 U9446 ( .A(n8191), .ZN(n7901) );
  NOR2_X4 U9447 ( .A1(n8193), .A2(n7901), .ZN(n8008) );
  OAI21_X4 U9448 ( .B1(n7906), .B2(n7905), .A(n7904), .ZN(n7907) );
  AOI21_X4 U9449 ( .B1(a[14]), .B2(b[20]), .A(n7907), .ZN(n8245) );
  NAND2_X2 U9450 ( .A1(a[14]), .A2(n7907), .ZN(n8243) );
  INV_X4 U9451 ( .A(n8243), .ZN(n7908) );
  NOR2_X4 U9452 ( .A1(n8245), .A2(n7908), .ZN(n8006) );
  INV_X4 U9453 ( .A(n7909), .ZN(n7911) );
  NOR2_X4 U9454 ( .A1(n7911), .A2(n7910), .ZN(n7913) );
  NAND2_X2 U9455 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  OAI21_X4 U9456 ( .B1(n7913), .B2(n8197), .A(n7912), .ZN(n8194) );
  XNOR2_X2 U9457 ( .A(n8195), .B(n8194), .ZN(n7915) );
  NAND2_X2 U9458 ( .A1(a[4]), .A2(net248517), .ZN(n8196) );
  INV_X4 U9459 ( .A(n8196), .ZN(n7914) );
  XNOR2_X2 U9460 ( .A(n7915), .B(n7914), .ZN(n8202) );
  NAND2_X2 U9461 ( .A1(a[5]), .A2(b[29]), .ZN(n7923) );
  INV_X4 U9462 ( .A(n7923), .ZN(n7921) );
  OAI21_X4 U9463 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n7922) );
  NAND2_X2 U9464 ( .A1(n7921), .A2(n7922), .ZN(n8201) );
  INV_X4 U9465 ( .A(n7922), .ZN(n7924) );
  NAND2_X2 U9466 ( .A1(n7924), .A2(n7923), .ZN(n8200) );
  NAND2_X2 U9467 ( .A1(n8201), .A2(n8200), .ZN(n7925) );
  XNOR2_X2 U9468 ( .A(n8202), .B(n7925), .ZN(n8206) );
  NAND2_X2 U9469 ( .A1(a[6]), .A2(net246880), .ZN(n7933) );
  INV_X4 U9470 ( .A(n7933), .ZN(n7931) );
  NOR2_X4 U9471 ( .A1(n7927), .A2(n7926), .ZN(n7930) );
  NAND2_X2 U9472 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  OAI21_X4 U9473 ( .B1(n7930), .B2(n7929), .A(n7928), .ZN(n7932) );
  NAND2_X2 U9474 ( .A1(n7931), .A2(n7932), .ZN(n8205) );
  INV_X4 U9475 ( .A(n7932), .ZN(n7934) );
  NAND2_X2 U9476 ( .A1(n7934), .A2(n7933), .ZN(n8204) );
  NAND2_X2 U9477 ( .A1(n8205), .A2(n8204), .ZN(n7935) );
  XNOR2_X2 U9478 ( .A(n8206), .B(n7935), .ZN(n8211) );
  NAND2_X2 U9479 ( .A1(a[7]), .A2(b[27]), .ZN(n7943) );
  INV_X4 U9480 ( .A(n7943), .ZN(n7941) );
  OAI21_X4 U9481 ( .B1(n7940), .B2(n7939), .A(n7938), .ZN(n7942) );
  NAND2_X2 U9482 ( .A1(n7941), .A2(n7942), .ZN(n8210) );
  INV_X4 U9483 ( .A(n7942), .ZN(n7944) );
  NAND2_X2 U9484 ( .A1(n7944), .A2(n7943), .ZN(n8209) );
  NAND2_X2 U9485 ( .A1(n8210), .A2(n8209), .ZN(n7945) );
  XNOR2_X2 U9486 ( .A(n8211), .B(n7945), .ZN(n8216) );
  NAND2_X2 U9487 ( .A1(a[8]), .A2(b[26]), .ZN(n7953) );
  INV_X4 U9488 ( .A(n7953), .ZN(n7951) );
  OAI21_X4 U9489 ( .B1(n7950), .B2(n7949), .A(n7948), .ZN(n7952) );
  NAND2_X2 U9490 ( .A1(n7951), .A2(n7952), .ZN(n8215) );
  INV_X4 U9491 ( .A(n7952), .ZN(n7954) );
  NAND2_X2 U9492 ( .A1(n7954), .A2(n7953), .ZN(n8214) );
  NAND2_X2 U9493 ( .A1(n8215), .A2(n8214), .ZN(n7955) );
  XNOR2_X2 U9494 ( .A(n8216), .B(n7955), .ZN(n8221) );
  NAND2_X2 U9495 ( .A1(a[9]), .A2(b[25]), .ZN(n7963) );
  INV_X4 U9496 ( .A(n7963), .ZN(n7961) );
  OAI21_X4 U9497 ( .B1(n7960), .B2(n7959), .A(n7958), .ZN(n7962) );
  NAND2_X2 U9498 ( .A1(n7961), .A2(n7962), .ZN(n8220) );
  INV_X4 U9499 ( .A(n7962), .ZN(n7964) );
  NAND2_X2 U9500 ( .A1(n7964), .A2(n7963), .ZN(n8219) );
  NAND2_X2 U9501 ( .A1(n8220), .A2(n8219), .ZN(n7965) );
  XNOR2_X2 U9502 ( .A(n8221), .B(n7965), .ZN(n8225) );
  NAND2_X2 U9503 ( .A1(a[10]), .A2(b[24]), .ZN(n7973) );
  INV_X4 U9504 ( .A(n7973), .ZN(n7971) );
  OAI21_X4 U9505 ( .B1(n7970), .B2(n7969), .A(n7968), .ZN(n7972) );
  NAND2_X2 U9506 ( .A1(n7971), .A2(n7972), .ZN(n8224) );
  INV_X4 U9507 ( .A(n7972), .ZN(n7974) );
  NAND2_X2 U9508 ( .A1(n7974), .A2(n7973), .ZN(n8223) );
  NAND2_X2 U9509 ( .A1(n8224), .A2(n8223), .ZN(n7975) );
  XNOR2_X2 U9510 ( .A(n8225), .B(n7975), .ZN(n8230) );
  NAND2_X2 U9511 ( .A1(a[11]), .A2(b[23]), .ZN(n7983) );
  INV_X4 U9512 ( .A(n7983), .ZN(n7981) );
  OAI21_X4 U9513 ( .B1(n7980), .B2(n7979), .A(n7978), .ZN(n7982) );
  NAND2_X2 U9514 ( .A1(n7981), .A2(n7982), .ZN(n8229) );
  INV_X4 U9515 ( .A(n7982), .ZN(n7984) );
  NAND2_X2 U9516 ( .A1(n7984), .A2(n7983), .ZN(n8228) );
  NAND2_X2 U9517 ( .A1(n8229), .A2(n8228), .ZN(n7985) );
  XNOR2_X2 U9518 ( .A(n8230), .B(n7985), .ZN(n8235) );
  NAND2_X2 U9519 ( .A1(a[12]), .A2(b[22]), .ZN(n7993) );
  INV_X4 U9520 ( .A(n7993), .ZN(n7991) );
  OAI21_X4 U9521 ( .B1(n7990), .B2(n7989), .A(n7988), .ZN(n7992) );
  NAND2_X2 U9522 ( .A1(n7991), .A2(n7992), .ZN(n8234) );
  INV_X4 U9523 ( .A(n7992), .ZN(n7994) );
  NAND2_X2 U9524 ( .A1(n7994), .A2(n7993), .ZN(n8233) );
  NAND2_X2 U9525 ( .A1(n8234), .A2(n8233), .ZN(n7995) );
  XNOR2_X2 U9526 ( .A(n8235), .B(n7995), .ZN(n8240) );
  NAND2_X2 U9527 ( .A1(a[13]), .A2(net246836), .ZN(n8003) );
  INV_X4 U9528 ( .A(n8003), .ZN(n8001) );
  NAND2_X2 U9529 ( .A1(n7997), .A2(n4423), .ZN(n7998) );
  NAND2_X2 U9530 ( .A1(n8001), .A2(n8002), .ZN(n8239) );
  INV_X4 U9531 ( .A(n8002), .ZN(n8004) );
  NAND2_X2 U9532 ( .A1(n8004), .A2(n8003), .ZN(n8238) );
  NAND2_X2 U9533 ( .A1(n8239), .A2(n8238), .ZN(n8005) );
  XNOR2_X2 U9534 ( .A(n8240), .B(n8005), .ZN(n8244) );
  XNOR2_X2 U9535 ( .A(n8006), .B(n8244), .ZN(n8007) );
  INV_X4 U9536 ( .A(n8007), .ZN(n8192) );
  XNOR2_X2 U9537 ( .A(n8008), .B(n8192), .ZN(n8188) );
  INV_X4 U9538 ( .A(n8188), .ZN(n8021) );
  NAND2_X2 U9539 ( .A1(n4578), .A2(b[18]), .ZN(n8017) );
  NAND3_X2 U9540 ( .A1(n8012), .A2(n8011), .A3(n8010), .ZN(n8013) );
  NAND3_X2 U9541 ( .A1(n8015), .A2(n8014), .A3(n8013), .ZN(n8016) );
  NAND2_X2 U9542 ( .A1(n8017), .A2(n8016), .ZN(n8187) );
  INV_X4 U9543 ( .A(n8016), .ZN(n8019) );
  INV_X4 U9544 ( .A(n8017), .ZN(n8018) );
  NAND2_X2 U9545 ( .A1(n8019), .A2(n8018), .ZN(n8189) );
  NAND2_X2 U9546 ( .A1(n8187), .A2(n8189), .ZN(n8020) );
  XNOR2_X2 U9547 ( .A(n8021), .B(n8020), .ZN(n8186) );
  INV_X4 U9548 ( .A(n8022), .ZN(n8023) );
  INV_X4 U9549 ( .A(n8183), .ZN(n8026) );
  XNOR2_X2 U9550 ( .A(n8026), .B(n8186), .ZN(n8027) );
  XNOR2_X2 U9551 ( .A(n8027), .B(n8182), .ZN(n8177) );
  INV_X4 U9552 ( .A(n8034), .ZN(n8028) );
  NOR2_X4 U9553 ( .A1(n8028), .A2(n4432), .ZN(n8030) );
  OAI21_X4 U9554 ( .B1(n8030), .B2(n8032), .A(n8029), .ZN(n8175) );
  NAND2_X2 U9555 ( .A1(n3979), .A2(n8175), .ZN(n8176) );
  OAI21_X4 U9556 ( .B1(n3979), .B2(n8175), .A(n8176), .ZN(n8172) );
  XNOR2_X2 U9557 ( .A(n8177), .B(n8172), .ZN(n8047) );
  NAND2_X2 U9558 ( .A1(b[15]), .A2(a[19]), .ZN(n8044) );
  INV_X4 U9559 ( .A(n8044), .ZN(n8042) );
  INV_X4 U9560 ( .A(n8031), .ZN(n8036) );
  XNOR2_X2 U9561 ( .A(n8033), .B(n8032), .ZN(n8035) );
  XNOR2_X2 U9562 ( .A(n8035), .B(n4451), .ZN(n8038) );
  NAND2_X2 U9563 ( .A1(n8036), .A2(n8038), .ZN(n8041) );
  NAND2_X2 U9564 ( .A1(n8036), .A2(n8037), .ZN(n8040) );
  NAND2_X2 U9565 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  INV_X4 U9566 ( .A(n8043), .ZN(n8045) );
  NAND2_X2 U9567 ( .A1(n8045), .A2(n8044), .ZN(n8173) );
  XNOR2_X2 U9568 ( .A(n8047), .B(n8046), .ZN(n8170) );
  XNOR2_X2 U9569 ( .A(n8050), .B(n8049), .ZN(n8051) );
  INV_X4 U9570 ( .A(n8051), .ZN(n8058) );
  INV_X4 U9571 ( .A(n8052), .ZN(n8056) );
  OAI21_X4 U9572 ( .B1(n8056), .B2(n8055), .A(n8054), .ZN(n8057) );
  NAND2_X2 U9573 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  OAI21_X4 U9574 ( .B1(n8061), .B2(n8060), .A(n8059), .ZN(n8064) );
  INV_X4 U9575 ( .A(n8064), .ZN(n8062) );
  NAND2_X2 U9576 ( .A1(a[20]), .A2(b[14]), .ZN(n8063) );
  NAND2_X2 U9577 ( .A1(n8062), .A2(n8063), .ZN(n8168) );
  INV_X4 U9578 ( .A(n8063), .ZN(n8065) );
  NAND2_X2 U9579 ( .A1(n8065), .A2(n8064), .ZN(n8169) );
  XNOR2_X2 U9580 ( .A(n8170), .B(n8066), .ZN(n8165) );
  NAND2_X2 U9581 ( .A1(b[13]), .A2(a[21]), .ZN(n8077) );
  INV_X4 U9582 ( .A(n8077), .ZN(n8075) );
  INV_X4 U9583 ( .A(n8067), .ZN(n8070) );
  NAND2_X2 U9584 ( .A1(n8075), .A2(n8076), .ZN(n8164) );
  INV_X4 U9585 ( .A(n8076), .ZN(n8078) );
  NAND2_X2 U9586 ( .A1(n8078), .A2(n8077), .ZN(n8163) );
  NAND2_X2 U9587 ( .A1(n8164), .A2(n8163), .ZN(n8079) );
  XNOR2_X2 U9588 ( .A(n8165), .B(n8079), .ZN(n8158) );
  INV_X4 U9589 ( .A(n8158), .ZN(n8144) );
  XNOR2_X2 U9590 ( .A(n8144), .B(n8145), .ZN(n8155) );
  NAND2_X2 U9591 ( .A1(b[11]), .A2(a[23]), .ZN(n8093) );
  INV_X4 U9592 ( .A(n8093), .ZN(n8091) );
  OAI21_X4 U9593 ( .B1(n8090), .B2(n3912), .A(n8089), .ZN(n8092) );
  NAND2_X2 U9594 ( .A1(n8091), .A2(n8092), .ZN(n8538) );
  INV_X4 U9595 ( .A(n8092), .ZN(n8094) );
  XNOR2_X2 U9596 ( .A(n8155), .B(n8268), .ZN(n8151) );
  INV_X4 U9597 ( .A(n8095), .ZN(n8099) );
  OAI21_X4 U9598 ( .B1(n8098), .B2(n8099), .A(n8097), .ZN(n8100) );
  NAND2_X2 U9599 ( .A1(a[24]), .A2(n8100), .ZN(net241493) );
  AOI21_X4 U9600 ( .B1(a[24]), .B2(b[10]), .A(n8100), .ZN(net241746) );
  XNOR2_X2 U9601 ( .A(n8151), .B(net241832), .ZN(n8102) );
  NAND2_X2 U9602 ( .A1(b[9]), .A2(net246760), .ZN(net241754) );
  INV_X4 U9603 ( .A(net241754), .ZN(net241749) );
  INV_X4 U9604 ( .A(net241760), .ZN(net241829) );
  NAND2_X2 U9605 ( .A1(net241830), .A2(net248509), .ZN(net241824) );
  INV_X4 U9606 ( .A(net241756), .ZN(net241827) );
  NAND2_X2 U9607 ( .A1(n8101), .A2(net241756), .ZN(net241596) );
  XNOR2_X2 U9608 ( .A(n8102), .B(net241821), .ZN(n8258) );
  XNOR2_X2 U9609 ( .A(net241581), .B(net241044), .ZN(n8103) );
  XNOR2_X2 U9610 ( .A(n4026), .B(n8103), .ZN(net241563) );
  NAND3_X4 U9611 ( .A1(n8104), .A2(a[31]), .A3(b[4]), .ZN(n8279) );
  XNOR2_X2 U9612 ( .A(n4057), .B(n8105), .ZN(n8280) );
  NAND2_X2 U9613 ( .A1(net240913), .A2(n8281), .ZN(n8108) );
  NAND2_X2 U9614 ( .A1(n8108), .A2(n4550), .ZN(n8129) );
  AOI22_X2 U9615 ( .A1(n8841), .A2(n8110), .B1(n8842), .B2(n8109), .ZN(n8127)
         );
  NAND2_X2 U9616 ( .A1(n8111), .A2(n4565), .ZN(n8114) );
  INV_X4 U9617 ( .A(n8112), .ZN(n8113) );
  OAI211_X2 U9618 ( .C1(n1323), .C2(n8115), .A(n8114), .B(n8113), .ZN(n8309)
         );
  NAND2_X2 U9619 ( .A1(n4558), .A2(n8797), .ZN(n8122) );
  AOI22_X2 U9620 ( .A1(net247082), .A2(a[19]), .B1(n8834), .B2(net246772), 
        .ZN(n8116) );
  OAI211_X2 U9621 ( .C1(net246958), .C2(n8289), .A(n8117), .B(n8116), .ZN(
        n8794) );
  NAND2_X2 U9622 ( .A1(n3977), .A2(n8794), .ZN(n8121) );
  NAND2_X2 U9623 ( .A1(n4562), .A2(n8118), .ZN(n8120) );
  NAND2_X2 U9624 ( .A1(n4555), .A2(n8795), .ZN(n8119) );
  NAND4_X2 U9625 ( .A1(n8122), .A2(n8121), .A3(n8120), .A4(n8119), .ZN(n8310)
         );
  INV_X4 U9626 ( .A(n8310), .ZN(n8123) );
  NAND2_X2 U9627 ( .A1(n8132), .A2(n8130), .ZN(n8135) );
  INV_X4 U9628 ( .A(n8131), .ZN(n8134) );
  INV_X4 U9629 ( .A(n8132), .ZN(n8133) );
  AOI22_X2 U9630 ( .A1(n8135), .A2(n8134), .B1(n8133), .B2(a[4]), .ZN(n8290)
         );
  XNOR2_X2 U9631 ( .A(net246924), .B(b[3]), .ZN(n8288) );
  XNOR2_X2 U9632 ( .A(a[3]), .B(n8288), .ZN(n8136) );
  XNOR2_X2 U9633 ( .A(n8290), .B(n8136), .ZN(n8140) );
  NAND2_X2 U9634 ( .A1(n8784), .A2(n8137), .ZN(n8138) );
  AOI21_X2 U9635 ( .B1(n4552), .B2(n8140), .A(n8139), .ZN(n8141) );
  OAI211_X2 U9636 ( .C1(n8143), .C2(n8281), .A(n8142), .B(n8141), .ZN(out[3])
         );
  XNOR2_X2 U9637 ( .A(n8144), .B(n8145), .ZN(n8539) );
  XNOR2_X2 U9638 ( .A(n4407), .B(n8268), .ZN(net241492) );
  NAND2_X2 U9639 ( .A1(n8146), .A2(net241756), .ZN(n8149) );
  INV_X4 U9640 ( .A(n8149), .ZN(n8147) );
  NAND2_X2 U9641 ( .A1(n8147), .A2(net241754), .ZN(n8148) );
  NAND2_X2 U9642 ( .A1(net241749), .A2(n8149), .ZN(n8327) );
  XNOR2_X2 U9643 ( .A(n3981), .B(n8150), .ZN(net241628) );
  NAND2_X2 U9644 ( .A1(a[23]), .A2(b[10]), .ZN(n8341) );
  INV_X4 U9645 ( .A(n8341), .ZN(n8153) );
  XNOR2_X2 U9646 ( .A(n8153), .B(n8152), .ZN(n8257) );
  INV_X4 U9647 ( .A(n8154), .ZN(n8540) );
  INV_X4 U9648 ( .A(n8156), .ZN(n8159) );
  OAI21_X4 U9649 ( .B1(n8159), .B2(n4399), .A(n8157), .ZN(n8535) );
  NAND2_X2 U9650 ( .A1(b[12]), .A2(a[21]), .ZN(n8534) );
  NAND2_X2 U9651 ( .A1(b[11]), .A2(a[22]), .ZN(n8544) );
  XNOR2_X2 U9652 ( .A(n8534), .B(n8544), .ZN(n8160) );
  XNOR2_X2 U9653 ( .A(n8535), .B(n8160), .ZN(n8161) );
  XNOR2_X2 U9654 ( .A(n8162), .B(n8161), .ZN(n8255) );
  INV_X4 U9655 ( .A(n8163), .ZN(n8166) );
  INV_X4 U9656 ( .A(n8517), .ZN(n8167) );
  NAND2_X2 U9657 ( .A1(b[13]), .A2(a[20]), .ZN(n8520) );
  XNOR2_X2 U9658 ( .A(n8167), .B(n8520), .ZN(n8253) );
  INV_X4 U9659 ( .A(n8168), .ZN(n8171) );
  NAND2_X2 U9660 ( .A1(a[19]), .A2(b[14]), .ZN(n8510) );
  XOR2_X2 U9661 ( .A(n8507), .B(n8510), .Z(n8252) );
  INV_X4 U9662 ( .A(n8173), .ZN(n8496) );
  NAND2_X2 U9663 ( .A1(b[15]), .A2(a[18]), .ZN(n8500) );
  XNOR2_X2 U9664 ( .A(n8174), .B(n8500), .ZN(n8251) );
  NAND2_X2 U9665 ( .A1(a[17]), .A2(b[16]), .ZN(n8490) );
  INV_X4 U9666 ( .A(n8490), .ZN(n8179) );
  NOR2_X4 U9667 ( .A1(n3979), .A2(n8175), .ZN(n8178) );
  OAI21_X4 U9668 ( .B1(n8178), .B2(n8177), .A(n8176), .ZN(n8487) );
  XNOR2_X2 U9669 ( .A(n8179), .B(n8487), .ZN(n8249) );
  NAND2_X2 U9670 ( .A1(b[17]), .A2(n4578), .ZN(n8480) );
  INV_X4 U9671 ( .A(n8182), .ZN(n8184) );
  NAND2_X2 U9672 ( .A1(n8184), .A2(n8183), .ZN(n8185) );
  OAI21_X4 U9673 ( .B1(n8186), .B2(n3948), .A(n8185), .ZN(n8477) );
  XOR2_X2 U9674 ( .A(n8480), .B(n8477), .Z(n8248) );
  NAND2_X2 U9675 ( .A1(n8188), .A2(n8187), .ZN(n8190) );
  NAND2_X2 U9676 ( .A1(n8190), .A2(n8189), .ZN(n8466) );
  NAND2_X2 U9677 ( .A1(a[15]), .A2(b[18]), .ZN(n8469) );
  XOR2_X2 U9678 ( .A(n8466), .B(n8469), .Z(n8247) );
  NAND2_X2 U9679 ( .A1(a[14]), .A2(b[19]), .ZN(n8458) );
  OAI21_X4 U9680 ( .B1(n8193), .B2(n8192), .A(n8191), .ZN(n8455) );
  XOR2_X2 U9681 ( .A(n8458), .B(n8455), .Z(n8246) );
  INV_X4 U9682 ( .A(n8194), .ZN(n8198) );
  NAND2_X2 U9683 ( .A1(a[3]), .A2(net248516), .ZN(n8348) );
  OAI21_X4 U9684 ( .B1(n8198), .B2(n3941), .A(n3974), .ZN(n8349) );
  XNOR2_X2 U9685 ( .A(n8348), .B(n8352), .ZN(n8199) );
  XNOR2_X2 U9686 ( .A(n8349), .B(n8199), .ZN(n8355) );
  INV_X4 U9687 ( .A(n8200), .ZN(n8203) );
  OAI21_X4 U9688 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8356) );
  NAND2_X2 U9689 ( .A1(a[4]), .A2(b[29]), .ZN(n8358) );
  INV_X4 U9690 ( .A(n8204), .ZN(n8207) );
  OAI21_X4 U9691 ( .B1(n8207), .B2(n8206), .A(n8205), .ZN(n8365) );
  XOR2_X2 U9692 ( .A(n8366), .B(n8365), .Z(n8208) );
  NAND2_X2 U9693 ( .A1(a[5]), .A2(net246880), .ZN(n8368) );
  XNOR2_X2 U9694 ( .A(n8208), .B(n8368), .ZN(n8375) );
  INV_X4 U9695 ( .A(n8209), .ZN(n8212) );
  OAI21_X4 U9696 ( .B1(n8212), .B2(n8211), .A(n8210), .ZN(n8376) );
  XOR2_X2 U9697 ( .A(n8375), .B(n8376), .Z(n8213) );
  NAND2_X2 U9698 ( .A1(a[6]), .A2(b[27]), .ZN(n8378) );
  XNOR2_X2 U9699 ( .A(n8213), .B(n8378), .ZN(n8386) );
  INV_X4 U9700 ( .A(n8214), .ZN(n8217) );
  OAI21_X4 U9701 ( .B1(n8217), .B2(n8216), .A(n8215), .ZN(n8385) );
  XOR2_X2 U9702 ( .A(n8386), .B(n8385), .Z(n8218) );
  NAND2_X2 U9703 ( .A1(a[7]), .A2(b[26]), .ZN(n8388) );
  XNOR2_X2 U9704 ( .A(n8218), .B(n8388), .ZN(n8395) );
  INV_X4 U9705 ( .A(n8219), .ZN(n8222) );
  OAI21_X4 U9706 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8396) );
  NAND2_X2 U9707 ( .A1(a[8]), .A2(b[25]), .ZN(n8398) );
  INV_X4 U9708 ( .A(n8223), .ZN(n8226) );
  OAI21_X4 U9709 ( .B1(n8226), .B2(n8225), .A(n8224), .ZN(n8405) );
  XOR2_X2 U9710 ( .A(n8406), .B(n8405), .Z(n8227) );
  NAND2_X2 U9711 ( .A1(a[9]), .A2(b[24]), .ZN(n8408) );
  XNOR2_X2 U9712 ( .A(n8227), .B(n8408), .ZN(n8415) );
  INV_X4 U9713 ( .A(n8228), .ZN(n8231) );
  OAI21_X4 U9714 ( .B1(n8231), .B2(n8230), .A(n8229), .ZN(n8416) );
  XOR2_X2 U9715 ( .A(n8415), .B(n8416), .Z(n8232) );
  NAND2_X2 U9716 ( .A1(a[10]), .A2(b[23]), .ZN(n8418) );
  XNOR2_X2 U9717 ( .A(n8232), .B(n8418), .ZN(n8426) );
  INV_X4 U9718 ( .A(n8233), .ZN(n8236) );
  OAI21_X4 U9719 ( .B1(n8236), .B2(n8235), .A(n8234), .ZN(n8425) );
  XOR2_X2 U9720 ( .A(n8426), .B(n8425), .Z(n8237) );
  NAND2_X2 U9721 ( .A1(a[11]), .A2(b[22]), .ZN(n8428) );
  XNOR2_X2 U9722 ( .A(n8237), .B(n8428), .ZN(n8435) );
  INV_X4 U9723 ( .A(n8238), .ZN(n8241) );
  OAI21_X4 U9724 ( .B1(n8241), .B2(n8240), .A(n8239), .ZN(n8436) );
  XOR2_X2 U9725 ( .A(n8435), .B(n8436), .Z(n8242) );
  NAND2_X2 U9726 ( .A1(a[12]), .A2(net246836), .ZN(n8438) );
  XNOR2_X2 U9727 ( .A(n8242), .B(n8438), .ZN(n8446) );
  OAI21_X4 U9728 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n8445) );
  NAND2_X2 U9729 ( .A1(a[13]), .A2(b[20]), .ZN(n8448) );
  XNOR2_X2 U9730 ( .A(n8246), .B(n8456), .ZN(n8467) );
  XNOR2_X2 U9731 ( .A(n8247), .B(n8467), .ZN(n8478) );
  XNOR2_X2 U9732 ( .A(n8248), .B(n8478), .ZN(n8488) );
  XNOR2_X2 U9733 ( .A(n8249), .B(n8488), .ZN(n8497) );
  INV_X4 U9734 ( .A(n8497), .ZN(n8250) );
  XNOR2_X2 U9735 ( .A(n8251), .B(n8250), .ZN(n8508) );
  XNOR2_X2 U9736 ( .A(n8252), .B(n8508), .ZN(n8518) );
  XNOR2_X2 U9737 ( .A(n8253), .B(n8518), .ZN(n8536) );
  XNOR2_X2 U9738 ( .A(n8255), .B(n8254), .ZN(n8337) );
  INV_X4 U9739 ( .A(n8337), .ZN(n8256) );
  XNOR2_X2 U9740 ( .A(n8257), .B(n8256), .ZN(net241503) );
  INV_X4 U9741 ( .A(n8266), .ZN(n8264) );
  NAND2_X2 U9742 ( .A1(n8259), .A2(net241625), .ZN(n8263) );
  INV_X4 U9743 ( .A(n8269), .ZN(n8260) );
  NAND2_X2 U9744 ( .A1(n8260), .A2(net241625), .ZN(n8261) );
  INV_X4 U9745 ( .A(n8265), .ZN(n8267) );
  INV_X4 U9746 ( .A(n8268), .ZN(n8270) );
  XNOR2_X2 U9747 ( .A(n8270), .B(n8269), .ZN(n8272) );
  XNOR2_X2 U9748 ( .A(n8272), .B(n8271), .ZN(net241597) );
  XNOR2_X2 U9749 ( .A(net241581), .B(net241044), .ZN(net241014) );
  OAI21_X4 U9750 ( .B1(n8275), .B2(n8274), .A(net241579), .ZN(net241013) );
  INV_X4 U9751 ( .A(n8278), .ZN(n8277) );
  NAND2_X2 U9752 ( .A1(n8277), .A2(n8276), .ZN(net241565) );
  NAND2_X2 U9753 ( .A1(b[4]), .A2(net246788), .ZN(net241566) );
  INV_X4 U9754 ( .A(net241566), .ZN(net241568) );
  NAND2_X2 U9755 ( .A1(n8279), .A2(n8278), .ZN(net241567) );
  XNOR2_X2 U9756 ( .A(net240961), .B(net241561), .ZN(n8770) );
  NAND2_X2 U9757 ( .A1(b[3]), .A2(a[30]), .ZN(n8766) );
  XNOR2_X2 U9758 ( .A(n8767), .B(n8766), .ZN(n8282) );
  XNOR2_X2 U9759 ( .A(n8770), .B(n8282), .ZN(n8772) );
  NAND2_X2 U9760 ( .A1(net240782), .A2(a[2]), .ZN(n8283) );
  NAND2_X2 U9761 ( .A1(net240913), .A2(net241554), .ZN(n8285) );
  NAND2_X2 U9762 ( .A1(n8285), .A2(n4550), .ZN(n8286) );
  NAND2_X2 U9763 ( .A1(n8784), .A2(n8287), .ZN(n8324) );
  XNOR2_X2 U9764 ( .A(net246924), .B(b[2]), .ZN(n8774) );
  XNOR2_X2 U9765 ( .A(a[2]), .B(n8774), .ZN(n8294) );
  INV_X4 U9766 ( .A(n8288), .ZN(n8292) );
  NAND2_X2 U9767 ( .A1(n8290), .A2(n8289), .ZN(n8291) );
  OAI21_X4 U9768 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8775) );
  XNOR2_X2 U9769 ( .A(n8294), .B(n8775), .ZN(n8322) );
  INV_X4 U9770 ( .A(n8295), .ZN(n8297) );
  NOR2_X4 U9771 ( .A1(n8297), .A2(n8296), .ZN(n8302) );
  NAND2_X2 U9772 ( .A1(n8302), .A2(n8301), .ZN(n8304) );
  MUX2_X2 U9773 ( .A(n8304), .B(n8303), .S(b[29]), .Z(n8839) );
  INV_X4 U9774 ( .A(n8839), .ZN(n8308) );
  NAND2_X2 U9775 ( .A1(n4555), .A2(n8831), .ZN(n8307) );
  NAND2_X2 U9776 ( .A1(n4561), .A2(n8305), .ZN(n8306) );
  OAI211_X2 U9777 ( .C1(net248517), .C2(n8308), .A(n8307), .B(n8306), .ZN(
        n8788) );
  INV_X4 U9778 ( .A(n8309), .ZN(n8313) );
  NAND2_X2 U9779 ( .A1(n8841), .A2(n8310), .ZN(n8311) );
  MUX2_X2 U9780 ( .A(n8845), .B(n8314), .S(n4564), .Z(n8802) );
  INV_X4 U9781 ( .A(n8802), .ZN(n8315) );
  AOI211_X2 U9782 ( .C1(n8318), .C2(n8788), .A(n8317), .B(n8316), .ZN(n8320)
         );
  NAND2_X2 U9783 ( .A1(n4267), .A2(a[2]), .ZN(n8319) );
  AOI21_X2 U9784 ( .B1(n4552), .B2(n8322), .A(n8321), .ZN(n8323) );
  NAND4_X2 U9785 ( .A1(n8326), .A2(n8325), .A3(n8324), .A4(n8323), .ZN(out[2])
         );
  NAND2_X2 U9786 ( .A1(b[9]), .A2(a[23]), .ZN(n8334) );
  INV_X4 U9787 ( .A(n8334), .ZN(n8332) );
  NAND2_X2 U9788 ( .A1(n8331), .A2(n8330), .ZN(n8333) );
  NAND2_X2 U9789 ( .A1(n8332), .A2(n8333), .ZN(n8557) );
  INV_X4 U9790 ( .A(n8333), .ZN(n8335) );
  NAND2_X2 U9791 ( .A1(n8335), .A2(n8334), .ZN(n8556) );
  NAND2_X2 U9792 ( .A1(n8557), .A2(n8556), .ZN(n8336) );
  INV_X4 U9793 ( .A(n8336), .ZN(n8757) );
  NAND2_X2 U9794 ( .A1(a[22]), .A2(b[10]), .ZN(n8345) );
  INV_X4 U9795 ( .A(n8345), .ZN(n8343) );
  INV_X4 U9796 ( .A(n4456), .ZN(n8339) );
  NOR2_X4 U9797 ( .A1(n8339), .A2(n8338), .ZN(n8342) );
  NAND2_X2 U9798 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  OAI21_X4 U9799 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8344) );
  NAND2_X2 U9800 ( .A1(n8343), .A2(n8344), .ZN(n8561) );
  INV_X4 U9801 ( .A(n8344), .ZN(n8346) );
  NAND2_X2 U9802 ( .A1(a[1]), .A2(net249231), .ZN(n8634) );
  INV_X4 U9803 ( .A(n8348), .ZN(n8350) );
  NOR2_X4 U9804 ( .A1(n8350), .A2(n8349), .ZN(n8353) );
  NAND2_X2 U9805 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  OAI21_X4 U9806 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8632) );
  XNOR2_X2 U9807 ( .A(n8634), .B(n8632), .ZN(n8354) );
  XNOR2_X2 U9808 ( .A(n3975), .B(n8354), .ZN(n8630) );
  NAND2_X2 U9809 ( .A1(a[3]), .A2(b[29]), .ZN(n8362) );
  INV_X4 U9810 ( .A(n8362), .ZN(n8360) );
  NOR2_X4 U9811 ( .A1(n8355), .A2(n8356), .ZN(n8359) );
  NAND2_X2 U9812 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  OAI21_X4 U9813 ( .B1(n8359), .B2(n8358), .A(n8357), .ZN(n8361) );
  NAND2_X2 U9814 ( .A1(n8360), .A2(n8361), .ZN(n8629) );
  INV_X4 U9815 ( .A(n8361), .ZN(n8363) );
  NAND2_X2 U9816 ( .A1(n8363), .A2(n8362), .ZN(n8628) );
  NAND2_X2 U9817 ( .A1(n8629), .A2(n8628), .ZN(n8364) );
  XNOR2_X2 U9818 ( .A(n8630), .B(n8364), .ZN(n8626) );
  NAND2_X2 U9819 ( .A1(a[4]), .A2(net246880), .ZN(n8372) );
  INV_X4 U9820 ( .A(n8372), .ZN(n8370) );
  NOR2_X4 U9821 ( .A1(n8366), .A2(n8365), .ZN(n8369) );
  NAND2_X2 U9822 ( .A1(n8366), .A2(n8365), .ZN(n8367) );
  OAI21_X4 U9823 ( .B1(n8369), .B2(n8368), .A(n8367), .ZN(n8371) );
  NAND2_X2 U9824 ( .A1(n8370), .A2(n8371), .ZN(n8625) );
  INV_X4 U9825 ( .A(n8371), .ZN(n8373) );
  NAND2_X2 U9826 ( .A1(n8373), .A2(n8372), .ZN(n8624) );
  NAND2_X2 U9827 ( .A1(n8625), .A2(n8624), .ZN(n8374) );
  XNOR2_X2 U9828 ( .A(n8626), .B(n8374), .ZN(n8622) );
  NAND2_X2 U9829 ( .A1(a[5]), .A2(b[27]), .ZN(n8382) );
  INV_X4 U9830 ( .A(n8382), .ZN(n8380) );
  NOR2_X4 U9831 ( .A1(n8375), .A2(n8376), .ZN(n8379) );
  NAND2_X2 U9832 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  OAI21_X4 U9833 ( .B1(n8379), .B2(n8378), .A(n8377), .ZN(n8381) );
  NAND2_X2 U9834 ( .A1(n8380), .A2(n8381), .ZN(n8621) );
  INV_X4 U9835 ( .A(n8381), .ZN(n8383) );
  NAND2_X2 U9836 ( .A1(n8383), .A2(n8382), .ZN(n8620) );
  NAND2_X2 U9837 ( .A1(n8621), .A2(n8620), .ZN(n8384) );
  XNOR2_X2 U9838 ( .A(n8622), .B(n8384), .ZN(n8618) );
  NAND2_X2 U9839 ( .A1(a[6]), .A2(b[26]), .ZN(n8392) );
  INV_X4 U9840 ( .A(n8392), .ZN(n8390) );
  NAND2_X2 U9841 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  OAI21_X4 U9842 ( .B1(n8389), .B2(n8388), .A(n8387), .ZN(n8391) );
  NAND2_X2 U9843 ( .A1(n8390), .A2(n8391), .ZN(n8617) );
  INV_X4 U9844 ( .A(n8391), .ZN(n8393) );
  NAND2_X2 U9845 ( .A1(n8393), .A2(n8392), .ZN(n8616) );
  NAND2_X2 U9846 ( .A1(n8617), .A2(n8616), .ZN(n8394) );
  XNOR2_X2 U9847 ( .A(n8618), .B(n8394), .ZN(n8614) );
  NAND2_X2 U9848 ( .A1(a[7]), .A2(b[25]), .ZN(n8402) );
  INV_X4 U9849 ( .A(n8402), .ZN(n8400) );
  NOR2_X4 U9850 ( .A1(n8395), .A2(n8396), .ZN(n8399) );
  NAND2_X2 U9851 ( .A1(n8396), .A2(n8395), .ZN(n8397) );
  OAI21_X4 U9852 ( .B1(n8399), .B2(n8398), .A(n8397), .ZN(n8401) );
  NAND2_X2 U9853 ( .A1(n8400), .A2(n8401), .ZN(n8613) );
  INV_X4 U9854 ( .A(n8401), .ZN(n8403) );
  NAND2_X2 U9855 ( .A1(n8403), .A2(n8402), .ZN(n8612) );
  NAND2_X2 U9856 ( .A1(n8613), .A2(n8612), .ZN(n8404) );
  XNOR2_X2 U9857 ( .A(n8614), .B(n8404), .ZN(n8610) );
  NAND2_X2 U9858 ( .A1(a[8]), .A2(b[24]), .ZN(n8412) );
  INV_X4 U9859 ( .A(n8412), .ZN(n8410) );
  NOR2_X4 U9860 ( .A1(n8406), .A2(n8405), .ZN(n8409) );
  NAND2_X2 U9861 ( .A1(n8406), .A2(n8405), .ZN(n8407) );
  OAI21_X4 U9862 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(n8411) );
  NAND2_X2 U9863 ( .A1(n8410), .A2(n8411), .ZN(n8609) );
  INV_X4 U9864 ( .A(n8411), .ZN(n8413) );
  NAND2_X2 U9865 ( .A1(n8413), .A2(n8412), .ZN(n8608) );
  NAND2_X2 U9866 ( .A1(n8609), .A2(n8608), .ZN(n8414) );
  XNOR2_X2 U9867 ( .A(n8610), .B(n8414), .ZN(n8606) );
  NAND2_X2 U9868 ( .A1(a[9]), .A2(b[23]), .ZN(n8422) );
  INV_X4 U9869 ( .A(n8422), .ZN(n8420) );
  NOR2_X4 U9870 ( .A1(n8415), .A2(n8416), .ZN(n8419) );
  NAND2_X2 U9871 ( .A1(n8416), .A2(n8415), .ZN(n8417) );
  OAI21_X4 U9872 ( .B1(n8419), .B2(n8418), .A(n8417), .ZN(n8421) );
  NAND2_X2 U9873 ( .A1(n8420), .A2(n8421), .ZN(n8605) );
  INV_X4 U9874 ( .A(n8421), .ZN(n8423) );
  NAND2_X2 U9875 ( .A1(n8423), .A2(n8422), .ZN(n8604) );
  NAND2_X2 U9876 ( .A1(n8605), .A2(n8604), .ZN(n8424) );
  XNOR2_X2 U9877 ( .A(n8606), .B(n8424), .ZN(n8602) );
  NAND2_X2 U9878 ( .A1(a[10]), .A2(b[22]), .ZN(n8432) );
  INV_X4 U9879 ( .A(n8432), .ZN(n8430) );
  OAI21_X4 U9880 ( .B1(n8429), .B2(n8428), .A(n8427), .ZN(n8431) );
  NAND2_X2 U9881 ( .A1(n8430), .A2(n8431), .ZN(n8601) );
  INV_X4 U9882 ( .A(n8431), .ZN(n8433) );
  NAND2_X2 U9883 ( .A1(n8433), .A2(n8432), .ZN(n8600) );
  NAND2_X2 U9884 ( .A1(n8601), .A2(n8600), .ZN(n8434) );
  XNOR2_X2 U9885 ( .A(n8602), .B(n8434), .ZN(n8598) );
  NAND2_X2 U9886 ( .A1(a[11]), .A2(net246836), .ZN(n8442) );
  INV_X4 U9887 ( .A(n8442), .ZN(n8440) );
  NAND2_X2 U9888 ( .A1(n8440), .A2(n8441), .ZN(n8597) );
  INV_X4 U9889 ( .A(n8441), .ZN(n8443) );
  NAND2_X2 U9890 ( .A1(n8443), .A2(n8442), .ZN(n8596) );
  NAND2_X2 U9891 ( .A1(n8597), .A2(n8596), .ZN(n8444) );
  XNOR2_X2 U9892 ( .A(n8598), .B(n8444), .ZN(n8594) );
  NAND2_X2 U9893 ( .A1(a[12]), .A2(b[20]), .ZN(n8452) );
  INV_X4 U9894 ( .A(n8452), .ZN(n8450) );
  NOR2_X4 U9895 ( .A1(n8446), .A2(n8445), .ZN(n8449) );
  NAND2_X2 U9896 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  OAI21_X4 U9897 ( .B1(n8449), .B2(n8448), .A(n8447), .ZN(n8451) );
  NAND2_X2 U9898 ( .A1(n8450), .A2(n8451), .ZN(n8593) );
  INV_X4 U9899 ( .A(n8451), .ZN(n8453) );
  NAND2_X2 U9900 ( .A1(n8453), .A2(n8452), .ZN(n8592) );
  NAND2_X2 U9901 ( .A1(n8593), .A2(n8592), .ZN(n8454) );
  XNOR2_X2 U9902 ( .A(n8594), .B(n8454), .ZN(n8590) );
  INV_X4 U9903 ( .A(n8590), .ZN(n8465) );
  NAND2_X2 U9904 ( .A1(a[13]), .A2(b[19]), .ZN(n8462) );
  INV_X4 U9905 ( .A(n8462), .ZN(n8460) );
  NAND2_X2 U9906 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  OAI21_X4 U9907 ( .B1(n8459), .B2(n8458), .A(n8457), .ZN(n8461) );
  NAND2_X2 U9908 ( .A1(n8460), .A2(n8461), .ZN(n8589) );
  INV_X4 U9909 ( .A(n8461), .ZN(n8463) );
  NAND2_X2 U9910 ( .A1(n8463), .A2(n8462), .ZN(n8588) );
  NAND2_X2 U9911 ( .A1(n8589), .A2(n8588), .ZN(n8464) );
  XNOR2_X2 U9912 ( .A(n8465), .B(n8464), .ZN(n8587) );
  INV_X4 U9913 ( .A(n8587), .ZN(n8476) );
  NAND2_X2 U9914 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  OAI21_X4 U9915 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8473) );
  INV_X4 U9916 ( .A(n8473), .ZN(n8471) );
  NAND2_X2 U9917 ( .A1(a[14]), .A2(b[18]), .ZN(n8472) );
  NAND2_X2 U9918 ( .A1(n8471), .A2(n8472), .ZN(n8586) );
  INV_X4 U9919 ( .A(n8472), .ZN(n8474) );
  NAND2_X2 U9920 ( .A1(n8474), .A2(n8473), .ZN(n8584) );
  NAND2_X2 U9921 ( .A1(n8586), .A2(n8584), .ZN(n8475) );
  XNOR2_X2 U9922 ( .A(n8476), .B(n8475), .ZN(n8724) );
  NAND2_X2 U9923 ( .A1(b[17]), .A2(a[15]), .ZN(n8484) );
  INV_X4 U9924 ( .A(n8484), .ZN(n8482) );
  NAND2_X2 U9925 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  OAI21_X4 U9926 ( .B1(n8481), .B2(n8480), .A(n8479), .ZN(n8483) );
  NAND2_X2 U9927 ( .A1(n8482), .A2(n8483), .ZN(n8723) );
  INV_X4 U9928 ( .A(n8483), .ZN(n8485) );
  NAND2_X2 U9929 ( .A1(n8485), .A2(n8484), .ZN(n8722) );
  XNOR2_X2 U9930 ( .A(n8724), .B(n8486), .ZN(n8730) );
  NAND2_X2 U9931 ( .A1(n8488), .A2(n8487), .ZN(n8489) );
  OAI21_X4 U9932 ( .B1(n8491), .B2(n8490), .A(n8489), .ZN(n8492) );
  INV_X4 U9933 ( .A(n8492), .ZN(n8728) );
  XNOR2_X2 U9934 ( .A(n8730), .B(n8728), .ZN(n8493) );
  XNOR2_X2 U9935 ( .A(n8493), .B(n8729), .ZN(n8582) );
  NAND2_X2 U9936 ( .A1(b[15]), .A2(a[17]), .ZN(n8504) );
  INV_X4 U9937 ( .A(n8504), .ZN(n8502) );
  NAND2_X2 U9938 ( .A1(n8502), .A2(n8503), .ZN(n8581) );
  INV_X4 U9939 ( .A(n8503), .ZN(n8505) );
  NAND2_X2 U9940 ( .A1(n8505), .A2(n8504), .ZN(n8580) );
  NAND2_X2 U9941 ( .A1(n8581), .A2(n8580), .ZN(n8506) );
  XNOR2_X2 U9942 ( .A(n8582), .B(n8506), .ZN(n8578) );
  NAND2_X2 U9943 ( .A1(a[18]), .A2(b[14]), .ZN(n8514) );
  INV_X4 U9944 ( .A(n8514), .ZN(n8512) );
  NAND2_X2 U9945 ( .A1(n8512), .A2(n8513), .ZN(n8577) );
  INV_X4 U9946 ( .A(n8513), .ZN(n8515) );
  NAND2_X2 U9947 ( .A1(n8515), .A2(n8514), .ZN(n8576) );
  NAND2_X2 U9948 ( .A1(n8577), .A2(n8576), .ZN(n8516) );
  XNOR2_X2 U9949 ( .A(n8578), .B(n8516), .ZN(n8574) );
  NAND2_X2 U9950 ( .A1(b[13]), .A2(a[19]), .ZN(n8524) );
  INV_X4 U9951 ( .A(n8524), .ZN(n8522) );
  NAND2_X2 U9952 ( .A1(n8522), .A2(n8523), .ZN(n8573) );
  INV_X4 U9953 ( .A(n8523), .ZN(n8525) );
  NAND2_X2 U9954 ( .A1(n8525), .A2(n8524), .ZN(n8572) );
  NAND2_X2 U9955 ( .A1(n8573), .A2(n8572), .ZN(n8526) );
  XNOR2_X2 U9956 ( .A(n8574), .B(n8526), .ZN(n8570) );
  NAND2_X2 U9957 ( .A1(b[12]), .A2(a[20]), .ZN(n8531) );
  INV_X4 U9958 ( .A(n8531), .ZN(n8529) );
  NAND2_X2 U9959 ( .A1(n8536), .A2(n8535), .ZN(n8527) );
  OAI21_X4 U9960 ( .B1(n8528), .B2(n8534), .A(n8527), .ZN(n8530) );
  NAND2_X2 U9961 ( .A1(n8529), .A2(n8530), .ZN(n8569) );
  INV_X4 U9962 ( .A(n8530), .ZN(n8532) );
  NAND2_X2 U9963 ( .A1(n8532), .A2(n8531), .ZN(n8568) );
  NAND2_X2 U9964 ( .A1(n8569), .A2(n8568), .ZN(n8533) );
  XNOR2_X2 U9965 ( .A(n8570), .B(n8533), .ZN(n8566) );
  NAND2_X2 U9966 ( .A1(b[11]), .A2(a[21]), .ZN(n8548) );
  INV_X4 U9967 ( .A(n8548), .ZN(n8546) );
  XOR2_X2 U9968 ( .A(n8535), .B(n8534), .Z(n8537) );
  XNOR2_X2 U9969 ( .A(n8536), .B(n8537), .ZN(n8542) );
  NAND2_X2 U9970 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  OAI21_X4 U9971 ( .B1(n8545), .B2(n8544), .A(n8543), .ZN(n8547) );
  NAND2_X2 U9972 ( .A1(n8546), .A2(n8547), .ZN(n8565) );
  INV_X4 U9973 ( .A(n8547), .ZN(n8549) );
  NAND2_X2 U9974 ( .A1(n8549), .A2(n8548), .ZN(n8564) );
  NAND2_X2 U9975 ( .A1(n8565), .A2(n8564), .ZN(n8550) );
  XNOR2_X2 U9976 ( .A(n8566), .B(n8550), .ZN(n8562) );
  XNOR2_X2 U9977 ( .A(n8755), .B(n8754), .ZN(n8558) );
  XNOR2_X2 U9978 ( .A(n8757), .B(n8558), .ZN(n8555) );
  INV_X4 U9979 ( .A(n8553), .ZN(n8551) );
  NAND2_X2 U9980 ( .A1(a[24]), .A2(b[8]), .ZN(n8552) );
  NAND2_X2 U9981 ( .A1(n8551), .A2(n8552), .ZN(n8752) );
  INV_X4 U9982 ( .A(n8552), .ZN(n8554) );
  AOI21_X4 U9983 ( .B1(n8555), .B2(n8752), .A(n3947), .ZN(n8750) );
  INV_X4 U9984 ( .A(n8556), .ZN(n8559) );
  INV_X4 U9985 ( .A(n8560), .ZN(n8563) );
  INV_X4 U9986 ( .A(n8564), .ZN(n8567) );
  INV_X4 U9987 ( .A(n8568), .ZN(n8571) );
  INV_X4 U9988 ( .A(n8572), .ZN(n8575) );
  INV_X4 U9989 ( .A(n8576), .ZN(n8579) );
  INV_X4 U9990 ( .A(n8580), .ZN(n8583) );
  INV_X4 U9991 ( .A(n8584), .ZN(n8585) );
  INV_X4 U9992 ( .A(n8588), .ZN(n8591) );
  INV_X4 U9993 ( .A(n8592), .ZN(n8595) );
  INV_X4 U9994 ( .A(n8596), .ZN(n8599) );
  INV_X4 U9995 ( .A(n8600), .ZN(n8603) );
  INV_X4 U9996 ( .A(n8604), .ZN(n8607) );
  INV_X4 U9997 ( .A(n8608), .ZN(n8611) );
  INV_X4 U9998 ( .A(n8612), .ZN(n8615) );
  INV_X4 U9999 ( .A(n8616), .ZN(n8619) );
  INV_X4 U10000 ( .A(n8620), .ZN(n8623) );
  INV_X4 U10001 ( .A(n8624), .ZN(n8627) );
  INV_X4 U10002 ( .A(n8628), .ZN(n8631) );
  NOR2_X4 U10003 ( .A1(n3975), .A2(n8632), .ZN(n8635) );
  NAND2_X2 U10004 ( .A1(n3975), .A2(n8632), .ZN(n8633) );
  OAI21_X4 U10005 ( .B1(n8635), .B2(n8634), .A(n8633), .ZN(n8697) );
  NAND2_X2 U10006 ( .A1(a[7]), .A2(b[24]), .ZN(n8637) );
  NAND2_X2 U10007 ( .A1(b[5]), .A2(net246766), .ZN(n8636) );
  XOR2_X2 U10008 ( .A(n8637), .B(n8636), .Z(n8641) );
  NAND2_X2 U10009 ( .A1(a[24]), .A2(b[7]), .ZN(n8639) );
  NAND2_X2 U10010 ( .A1(a[6]), .A2(b[25]), .ZN(n8638) );
  XNOR2_X2 U10011 ( .A(n8639), .B(n8638), .ZN(n8640) );
  XNOR2_X2 U10012 ( .A(n8641), .B(n8640), .ZN(n8649) );
  NAND2_X2 U10013 ( .A1(b[3]), .A2(a[28]), .ZN(n8643) );
  NAND2_X2 U10014 ( .A1(net246772), .A2(b[4]), .ZN(n8642) );
  XNOR2_X2 U10015 ( .A(n8643), .B(n8642), .ZN(n8647) );
  NAND2_X2 U10016 ( .A1(a[23]), .A2(b[8]), .ZN(n8645) );
  NAND2_X2 U10017 ( .A1(a[21]), .A2(b[10]), .ZN(n8644) );
  XNOR2_X2 U10018 ( .A(n8645), .B(n8644), .ZN(n8646) );
  XNOR2_X2 U10019 ( .A(n8647), .B(n8646), .ZN(n8648) );
  XNOR2_X2 U10020 ( .A(n8649), .B(n8648), .ZN(n8665) );
  NAND2_X2 U10021 ( .A1(b[6]), .A2(net246760), .ZN(n8651) );
  NAND2_X2 U10022 ( .A1(a[5]), .A2(b[26]), .ZN(n8650) );
  XOR2_X2 U10023 ( .A(n8651), .B(n8650), .Z(n8655) );
  NAND2_X2 U10024 ( .A1(a[4]), .A2(b[27]), .ZN(n8653) );
  NAND2_X2 U10025 ( .A1(net246788), .A2(b[2]), .ZN(n8652) );
  XNOR2_X2 U10026 ( .A(n8653), .B(n8652), .ZN(n8654) );
  XNOR2_X2 U10027 ( .A(n8655), .B(n8654), .ZN(n8663) );
  NAND2_X2 U10028 ( .A1(a[2]), .A2(b[29]), .ZN(n8657) );
  XNOR2_X2 U10029 ( .A(n8657), .B(n8656), .ZN(n8661) );
  NAND2_X2 U10030 ( .A1(a[0]), .A2(net246916), .ZN(n8659) );
  NAND2_X2 U10031 ( .A1(a[3]), .A2(net246880), .ZN(n8658) );
  XNOR2_X2 U10032 ( .A(n8659), .B(n8658), .ZN(n8660) );
  XNOR2_X2 U10033 ( .A(n8661), .B(n8660), .ZN(n8662) );
  XNOR2_X2 U10034 ( .A(n8663), .B(n8662), .ZN(n8664) );
  XNOR2_X2 U10035 ( .A(n8665), .B(n8664), .ZN(n8695) );
  NAND2_X2 U10036 ( .A1(a[10]), .A2(net246836), .ZN(n8667) );
  NAND2_X2 U10037 ( .A1(b[11]), .A2(a[20]), .ZN(n8666) );
  XOR2_X2 U10038 ( .A(n8667), .B(n8666), .Z(n8671) );
  NAND2_X2 U10039 ( .A1(b[13]), .A2(a[18]), .ZN(n8669) );
  NAND2_X2 U10040 ( .A1(b[12]), .A2(a[19]), .ZN(n8668) );
  XNOR2_X2 U10041 ( .A(n8669), .B(n8668), .ZN(n8670) );
  XNOR2_X2 U10042 ( .A(n8671), .B(n8670), .ZN(n8679) );
  NAND2_X2 U10043 ( .A1(b[17]), .A2(a[14]), .ZN(n8673) );
  NAND2_X2 U10044 ( .A1(a[15]), .A2(b[16]), .ZN(n8672) );
  XOR2_X2 U10045 ( .A(n8673), .B(n8672), .Z(n8677) );
  NAND2_X2 U10046 ( .A1(b[9]), .A2(a[22]), .ZN(n8675) );
  NAND2_X2 U10047 ( .A1(a[8]), .A2(b[23]), .ZN(n8674) );
  XNOR2_X2 U10048 ( .A(n8675), .B(n8674), .ZN(n8676) );
  XNOR2_X2 U10049 ( .A(n8677), .B(n8676), .ZN(n8678) );
  XNOR2_X2 U10050 ( .A(n8679), .B(n8678), .ZN(n8693) );
  NAND2_X2 U10051 ( .A1(b[15]), .A2(n4578), .ZN(n8681) );
  NAND2_X2 U10052 ( .A1(a[17]), .A2(b[14]), .ZN(n8680) );
  XNOR2_X2 U10053 ( .A(n8681), .B(n8680), .ZN(n8685) );
  NAND2_X2 U10054 ( .A1(a[9]), .A2(b[22]), .ZN(n8683) );
  NAND2_X2 U10055 ( .A1(a[12]), .A2(b[19]), .ZN(n8682) );
  XNOR2_X2 U10056 ( .A(n8683), .B(n8682), .ZN(n8684) );
  XNOR2_X2 U10057 ( .A(n8685), .B(n8684), .ZN(n8691) );
  NAND2_X2 U10058 ( .A1(a[13]), .A2(b[18]), .ZN(n8687) );
  NAND2_X2 U10059 ( .A1(a[11]), .A2(b[20]), .ZN(n8686) );
  XNOR2_X2 U10060 ( .A(n8687), .B(n8686), .ZN(n8689) );
  NAND2_X2 U10061 ( .A1(a[1]), .A2(net246902), .ZN(n8688) );
  XNOR2_X2 U10062 ( .A(n8689), .B(n8688), .ZN(n8690) );
  XNOR2_X2 U10063 ( .A(n8691), .B(n8690), .ZN(n8692) );
  XNOR2_X2 U10064 ( .A(n8693), .B(n8692), .ZN(n8694) );
  XNOR2_X2 U10065 ( .A(n8695), .B(n8694), .ZN(n8696) );
  XNOR2_X2 U10066 ( .A(n8697), .B(n8696), .ZN(n8698) );
  XNOR2_X2 U10067 ( .A(n8699), .B(n8698), .ZN(n8700) );
  XNOR2_X2 U10068 ( .A(n8701), .B(n8700), .ZN(n8702) );
  XNOR2_X2 U10069 ( .A(n8703), .B(n8702), .ZN(n8704) );
  XNOR2_X2 U10070 ( .A(n8705), .B(n8704), .ZN(n8706) );
  XNOR2_X2 U10071 ( .A(n8707), .B(n8706), .ZN(n8708) );
  XNOR2_X2 U10072 ( .A(n8709), .B(n8708), .ZN(n8710) );
  XNOR2_X2 U10073 ( .A(n8711), .B(n8710), .ZN(n8712) );
  XNOR2_X2 U10074 ( .A(n8713), .B(n8712), .ZN(n8714) );
  XNOR2_X2 U10075 ( .A(n8715), .B(n8714), .ZN(n8716) );
  XNOR2_X2 U10076 ( .A(n8717), .B(n8716), .ZN(n8718) );
  XNOR2_X2 U10077 ( .A(n8719), .B(n8718), .ZN(n8720) );
  XNOR2_X2 U10078 ( .A(n8721), .B(n8720), .ZN(n8727) );
  INV_X4 U10079 ( .A(n8722), .ZN(n8725) );
  XNOR2_X2 U10080 ( .A(n8727), .B(n8726), .ZN(n8734) );
  NOR2_X4 U10081 ( .A1(n8732), .A2(n8731), .ZN(n8733) );
  XNOR2_X2 U10082 ( .A(n8734), .B(n8733), .ZN(n8735) );
  XNOR2_X2 U10083 ( .A(n8736), .B(n8735), .ZN(n8737) );
  XNOR2_X2 U10084 ( .A(n8738), .B(n8737), .ZN(n8739) );
  XNOR2_X2 U10085 ( .A(n8740), .B(n8739), .ZN(n8741) );
  XNOR2_X2 U10086 ( .A(n8742), .B(n8741), .ZN(n8743) );
  XNOR2_X2 U10087 ( .A(n8744), .B(n8743), .ZN(n8745) );
  XNOR2_X2 U10088 ( .A(n8746), .B(n8745), .ZN(n8747) );
  XNOR2_X2 U10089 ( .A(n8748), .B(n8747), .ZN(n8749) );
  XNOR2_X2 U10090 ( .A(n8750), .B(n8749), .ZN(n8760) );
  INV_X4 U10091 ( .A(net241069), .ZN(net241065) );
  NAND2_X2 U10092 ( .A1(net241065), .A2(n8751), .ZN(net241064) );
  INV_X4 U10093 ( .A(net241050), .ZN(net241061) );
  INV_X4 U10094 ( .A(n8752), .ZN(n8753) );
  NOR2_X4 U10095 ( .A1(n8753), .A2(n3947), .ZN(net241052) );
  XNOR2_X2 U10096 ( .A(n8757), .B(n8756), .ZN(net241053) );
  XNOR2_X2 U10097 ( .A(net241053), .B(net241052), .ZN(net240997) );
  INV_X4 U10098 ( .A(n8758), .ZN(n8759) );
  NAND2_X2 U10099 ( .A1(n8759), .A2(net241050), .ZN(net240995) );
  XNOR2_X2 U10100 ( .A(net241047), .B(n8760), .ZN(net241026) );
  NAND3_X4 U10101 ( .A1(net241036), .A2(n8761), .A3(net241038), .ZN(net241031)
         );
  INV_X4 U10102 ( .A(net241032), .ZN(net241030) );
  XNOR2_X2 U10103 ( .A(net240989), .B(net240990), .ZN(n8762) );
  XNOR2_X2 U10104 ( .A(n8762), .B(net240988), .ZN(n8763) );
  INV_X4 U10105 ( .A(net240980), .ZN(net240982) );
  NAND2_X2 U10106 ( .A1(net240978), .A2(n8763), .ZN(n8764) );
  INV_X4 U10107 ( .A(n8766), .ZN(n8768) );
  OAI21_X4 U10108 ( .B1(n8771), .B2(n8770), .A(n8769), .ZN(net240951) );
  NAND2_X2 U10109 ( .A1(b[3]), .A2(net246788), .ZN(net240952) );
  XNOR2_X2 U10110 ( .A(net240927), .B(net240928), .ZN(net240783) );
  INV_X4 U10111 ( .A(net240762), .ZN(net240775) );
  AOI21_X4 U10112 ( .B1(net240910), .B2(n4550), .A(net240912), .ZN(net240772)
         );
  NAND2_X2 U10113 ( .A1(n8775), .A2(n8773), .ZN(n8778) );
  INV_X4 U10114 ( .A(n8774), .ZN(n8777) );
  INV_X4 U10115 ( .A(n8775), .ZN(n8776) );
  AOI22_X2 U10116 ( .A1(n8778), .A2(n8777), .B1(n8776), .B2(a[2]), .ZN(n8827)
         );
  XNOR2_X2 U10117 ( .A(net246926), .B(b[1]), .ZN(n8826) );
  XNOR2_X2 U10118 ( .A(a[1]), .B(n8826), .ZN(n8779) );
  XNOR2_X2 U10119 ( .A(n8827), .B(n8779), .ZN(n8780) );
  NAND2_X2 U10120 ( .A1(n4552), .A2(n8780), .ZN(n8782) );
  INV_X4 U10121 ( .A(n8782), .ZN(n8864) );
  NAND2_X2 U10122 ( .A1(net247002), .A2(a[1]), .ZN(n8863) );
  NAND2_X2 U10123 ( .A1(n8784), .A2(n8783), .ZN(n8861) );
  NAND2_X2 U10124 ( .A1(n8863), .A2(n8861), .ZN(n8785) );
  NOR4_X2 U10125 ( .A1(out[28]), .A2(out[29]), .A3(out[30]), .A4(n8785), .ZN(
        n8809) );
  INV_X4 U10126 ( .A(n8787), .ZN(n8807) );
  INV_X4 U10127 ( .A(n8788), .ZN(n8805) );
  INV_X4 U10128 ( .A(n8789), .ZN(n8790) );
  AOI21_X4 U10129 ( .B1(net246960), .B2(a[1]), .A(n8790), .ZN(n8791) );
  AOI21_X4 U10130 ( .B1(n4555), .B2(n8794), .A(n8793), .ZN(n8799) );
  AOI22_X2 U10131 ( .A1(n4561), .A2(n8797), .B1(n4557), .B2(n8795), .ZN(n8798)
         );
  NAND2_X2 U10132 ( .A1(n8799), .A2(n8798), .ZN(n8840) );
  INV_X4 U10133 ( .A(n8840), .ZN(n8800) );
  NOR2_X4 U10134 ( .A1(n8800), .A2(n4537), .ZN(n8801) );
  AOI21_X4 U10135 ( .B1(n8842), .B2(n8802), .A(n8801), .ZN(n8803) );
  OAI221_X2 U10136 ( .B1(n8807), .B2(n4535), .C1(n8805), .C2(n4539), .A(n8803), 
        .ZN(n8808) );
  NAND2_X2 U10137 ( .A1(n4549), .A2(n8808), .ZN(n8867) );
  NAND2_X2 U10138 ( .A1(n8809), .A2(n8867), .ZN(n8810) );
  INV_X4 U10139 ( .A(out[26]), .ZN(n8811) );
  NAND2_X2 U10140 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  NOR2_X4 U10141 ( .A1(out[25]), .A2(n8813), .ZN(n8815) );
  INV_X4 U10142 ( .A(out[24]), .ZN(n8814) );
  NAND2_X2 U10143 ( .A1(n8815), .A2(n8814), .ZN(n8816) );
  NOR2_X4 U10144 ( .A1(out[23]), .A2(n8816), .ZN(n8818) );
  INV_X4 U10145 ( .A(out[22]), .ZN(n8817) );
  NAND2_X2 U10146 ( .A1(n8818), .A2(n8817), .ZN(n8819) );
  NOR2_X4 U10147 ( .A1(out[21]), .A2(n8819), .ZN(n8821) );
  INV_X4 U10148 ( .A(out[20]), .ZN(n8820) );
  NAND2_X2 U10149 ( .A1(n8821), .A2(n8820), .ZN(n8822) );
  NOR3_X4 U10150 ( .A1(out[31]), .A2(out[19]), .A3(n8822), .ZN(n8824) );
  INV_X4 U10151 ( .A(out[18]), .ZN(n8823) );
  NAND2_X2 U10152 ( .A1(n8824), .A2(n8823), .ZN(n8825) );
  NOR3_X4 U10153 ( .A1(n8864), .A2(out[17]), .A3(n8825), .ZN(net240812) );
  INV_X4 U10154 ( .A(out[16]), .ZN(net240813) );
  NOR2_X4 U10155 ( .A1(n8829), .A2(n8828), .ZN(n8830) );
  FA_X1 U10156 ( .A(n8830), .B(n8851), .CI(net246932), .S(n8857) );
  NAND2_X2 U10157 ( .A1(net240782), .A2(n8845), .ZN(n8855) );
  INV_X4 U10158 ( .A(n8831), .ZN(n8833) );
  AOI22_X2 U10159 ( .A1(net247082), .A2(a[16]), .B1(n8834), .B2(a[24]), .ZN(
        n8835) );
  OAI211_X2 U10160 ( .C1(net246958), .C2(net240839), .A(n8836), .B(n8835), 
        .ZN(n8837) );
  AOI211_X2 U10161 ( .C1(net246902), .C2(n8839), .A(n8838), .B(n3998), .ZN(
        n8849) );
  NAND2_X2 U10162 ( .A1(n8841), .A2(n8840), .ZN(n8847) );
  NAND2_X2 U10163 ( .A1(n8842), .A2(n4565), .ZN(n8843) );
  OAI211_X2 U10164 ( .C1(n8849), .C2(n4537), .A(n8847), .B(n8846), .ZN(n8853)
         );
  AOI21_X2 U10165 ( .B1(n4548), .B2(n8853), .A(n8852), .ZN(n8854) );
  OAI211_X2 U10166 ( .C1(n8857), .C2(n8856), .A(n8855), .B(n8854), .ZN(
        net240814) );
  INV_X4 U10167 ( .A(net240814), .ZN(net240761) );
  NAND2_X2 U10168 ( .A1(net240782), .A2(a[1]), .ZN(n8858) );
  NAND2_X2 U10169 ( .A1(n8858), .A2(net247048), .ZN(n8859) );
  INV_X4 U10170 ( .A(n8861), .ZN(n8862) );
  INV_X4 U10171 ( .A(n8863), .ZN(n8865) );
  NAND4_X2 U10172 ( .A1(n8868), .A2(n8867), .A3(n8866), .A4(net240767), .ZN(
        out[1]) );
endmodule

