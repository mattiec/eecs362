module mult32bit(a, b, prod);
	parameter width = 32;
	
	input [width-1:0] a, b;
	output [width-1:0] prod;
	
	
	wire [width-1:0] c0, s0;
	
	fa add000(0, a[0]&b[0], 0, prod[0], c0[0]);
	fa add001(0, a[1]&b[0], c0[0], s0[1], c0[1]);
	fa add002(0, a[2]&b[0], c0[1], s0[2], c0[2]);
	fa add003(0, a[3]&b[0], c0[2], s0[3], c0[3]);
	fa add004(0, a[4]&b[0], c0[3], s0[4], c0[4]);
	fa add005(0, a[5]&b[0], c0[4], s0[5], c0[5]);
	fa add006(0, a[6]&b[0], c0[5], s0[6], c0[6]);
	fa add007(0, a[7]&b[0], c0[6], s0[7], c0[7]);
	fa add008(0, a[8]&b[0], c0[7], s0[8], c0[8]);
	fa add009(0, a[9]&b[0], c0[8], s0[9], c0[9]);
	fa add010(0, a[10]&b[0], c0[9], s0[10], c0[10]);
	fa add011(0, a[11]&b[0], c0[10], s0[11], c0[11]);
	fa add012(0, a[12]&b[0], c0[11], s0[12], c0[12]);
	fa add013(0, a[13]&b[0], c0[12], s0[13], c0[13]);
	fa add014(0, a[14]&b[0], c0[13], s0[14], c0[14]);
	fa add015(0, a[15]&b[0], c0[14], s0[15], c0[15]);
	fa add016(0, a[16]&b[0], c0[15], s0[16], c0[16]);
	fa add017(0, a[17]&b[0], c0[16], s0[17], c0[17]);
	fa add018(0, a[18]&b[0], c0[17], s0[18], c0[18]);
	fa add019(0, a[19]&b[0], c0[18], s0[19], c0[19]);
	fa add020(0, a[20]&b[0], c0[19], s0[20], c0[20]);
	fa add021(0, a[21]&b[0], c0[20], s0[21], c0[21]);
	fa add022(0, a[22]&b[0], c0[21], s0[22], c0[22]);
	fa add023(0, a[23]&b[0], c0[22], s0[23], c0[23]);
	fa add024(0, a[24]&b[0], c0[23], s0[24], c0[24]);
	fa add025(0, a[25]&b[0], c0[24], s0[25], c0[25]);
	fa add026(0, a[26]&b[0], c0[25], s0[26], c0[26]);
	fa add027(0, a[27]&b[0], c0[26], s0[27], c0[27]);
	fa add028(0, a[28]&b[0], c0[27], s0[28], c0[28]);
	fa add029(0, a[29]&b[0], c0[28], s0[29], c0[29]);
	fa add030(0, a[30]&b[0], c0[29], s0[30], c0[30]);
	fa add031(0, a[31]&b[0], c0[30], s0[31], c0[31]);

	
	wire [width-1:0] c1, s1;

	fa add100(s0[1], a[0]&b[1], 0, prod[1], c1[0]);
	fa add101(s0[2], a[1]&b[1], c1[0], s1[1], c1[1]);
	fa add102(s0[3], a[2]&b[1], c1[1], s1[2], c1[2]);
	fa add103(s0[4], a[3]&b[1], c1[2], s1[3], c1[3]);
	fa add104(s0[5], a[4]&b[1], c1[3], s1[4], c1[4]);
	fa add105(s0[6], a[5]&b[1], c1[4], s1[5], c1[5]);
	fa add106(s0[7], a[6]&b[1], c1[5], s1[6], c1[6]);
	fa add107(s0[8], a[7]&b[1], c1[6], s1[7], c1[7]);
	fa add108(s0[9], a[8]&b[1], c1[7], s1[8], c1[8]);
	fa add109(s0[10], a[9]&b[1], c1[8], s1[9], c1[9]);
	fa add110(s0[11], a[10]&b[1], c1[9], s1[10], c1[10]);
	fa add111(s0[12], a[11]&b[1], c1[10], s1[11], c1[11]);
	fa add112(s0[13], a[12]&b[1], c1[11], s1[12], c1[12]);
	fa add113(s0[14], a[13]&b[1], c1[12], s1[13], c1[13]);
	fa add114(s0[15], a[14]&b[1], c1[13], s1[14], c1[14]);
	fa add115(s0[16], a[15]&b[1], c1[14], s1[15], c1[15]);
	fa add116(s0[17], a[16]&b[1], c1[15], s1[16], c1[16]);
	fa add117(s0[18], a[17]&b[1], c1[16], s1[17], c1[17]);
	fa add118(s0[19], a[18]&b[1], c1[17], s1[18], c1[18]);
	fa add119(s0[20], a[19]&b[1], c1[18], s1[19], c1[19]);
	fa add120(s0[21], a[20]&b[1], c1[19], s1[20], c1[20]);
	fa add121(s0[22], a[21]&b[1], c1[20], s1[21], c1[21]);
	fa add122(s0[23], a[22]&b[1], c1[21], s1[22], c1[22]);
	fa add123(s0[24], a[23]&b[1], c1[22], s1[23], c1[23]);
	fa add124(s0[25], a[24]&b[1], c1[23], s1[24], c1[24]);
	fa add125(s0[26], a[25]&b[1], c1[24], s1[25], c1[25]);
	fa add126(s0[27], a[26]&b[1], c1[25], s1[26], c1[26]);
	fa add127(s0[28], a[27]&b[1], c1[26], s1[27], c1[27]);
	fa add128(s0[29], a[28]&b[1], c1[27], s1[28], c1[28]);
	fa add129(s0[30], a[29]&b[1], c1[28], s1[29], c1[29]);
	fa add130(s0[31], a[30]&b[1], c1[29], s1[30], c1[30]);
	fa add131(0, a[31]&b[1], c1[30], s1[31], c1[31]);

	
	wire [width-1:0] c2, s2;

	fa add200(s1[1], a[0]&b[2], 0, prod[2], c2[0]);
	fa add201(s1[2], a[1]&b[2], c2[0], s2[1], c2[1]);
	fa add202(s1[3], a[2]&b[2], c2[1], s2[2], c2[2]);
	fa add203(s1[4], a[3]&b[2], c2[2], s2[3], c2[3]);
	fa add204(s1[5], a[4]&b[2], c2[3], s2[4], c2[4]);
	fa add205(s1[6], a[5]&b[2], c2[4], s2[5], c2[5]);
	fa add206(s1[7], a[6]&b[2], c2[5], s2[6], c2[6]);
	fa add207(s1[8], a[7]&b[2], c2[6], s2[7], c2[7]);
	fa add208(s1[9], a[8]&b[2], c2[7], s2[8], c2[8]);
	fa add209(s1[10], a[9]&b[2], c2[8], s2[9], c2[9]);
	fa add210(s1[11], a[10]&b[2], c2[9], s2[10], c2[10]);
	fa add211(s1[12], a[11]&b[2], c2[10], s2[11], c2[11]);
	fa add212(s1[13], a[12]&b[2], c2[11], s2[12], c2[12]);
	fa add213(s1[14], a[13]&b[2], c2[12], s2[13], c2[13]);
	fa add214(s1[15], a[14]&b[2], c2[13], s2[14], c2[14]);
	fa add215(s1[16], a[15]&b[2], c2[14], s2[15], c2[15]);
	fa add216(s1[17], a[16]&b[2], c2[15], s2[16], c2[16]);
	fa add217(s1[18], a[17]&b[2], c2[16], s2[17], c2[17]);
	fa add218(s1[19], a[18]&b[2], c2[17], s2[18], c2[18]);
	fa add219(s1[20], a[19]&b[2], c2[18], s2[19], c2[19]);
	fa add220(s1[21], a[20]&b[2], c2[19], s2[20], c2[20]);
	fa add221(s1[22], a[21]&b[2], c2[20], s2[21], c2[21]);
	fa add222(s1[23], a[22]&b[2], c2[21], s2[22], c2[22]);
	fa add223(s1[24], a[23]&b[2], c2[22], s2[23], c2[23]);
	fa add224(s1[25], a[24]&b[2], c2[23], s2[24], c2[24]);
	fa add225(s1[26], a[25]&b[2], c2[24], s2[25], c2[25]);
	fa add226(s1[27], a[26]&b[2], c2[25], s2[26], c2[26]);
	fa add227(s1[28], a[27]&b[2], c2[26], s2[27], c2[27]);
	fa add228(s1[29], a[28]&b[2], c2[27], s2[28], c2[28]);
	fa add229(s1[30], a[29]&b[2], c2[28], s2[29], c2[29]);
	fa add230(s1[31], a[30]&b[2], c2[29], s2[30], c2[30]);
	fa add231(0, a[31]&b[2], c2[30], s2[31], c2[31]);
	
	
	wire [width-1:0] c3, s3;

	fa add300(s2[1], a[0]&b[3], 0, prod[3], c3[0]);
	fa add301(s2[2], a[1]&b[3], c3[0], s3[1], c3[1]);
	fa add302(s2[3], a[2]&b[3], c3[1], s3[2], c3[2]);
	fa add303(s2[4], a[3]&b[3], c3[2], s3[3], c3[3]);
	fa add304(s2[5], a[4]&b[3], c3[3], s3[4], c3[4]);
	fa add305(s2[6], a[5]&b[3], c3[4], s3[5], c3[5]);
	fa add306(s2[7], a[6]&b[3], c3[5], s3[6], c3[6]);
	fa add307(s2[8], a[7]&b[3], c3[6], s3[7], c3[7]);
	fa add308(s2[9], a[8]&b[3], c3[7], s3[8], c3[8]);
	fa add309(s2[10], a[9]&b[3], c3[8], s3[9], c3[9]);
	fa add310(s2[11], a[10]&b[3], c3[9], s3[10], c3[10]);
	fa add311(s2[12], a[11]&b[3], c3[10], s3[11], c3[11]);
	fa add312(s2[13], a[12]&b[3], c3[11], s3[12], c3[12]);
	fa add313(s2[14], a[13]&b[3], c3[12], s3[13], c3[13]);
	fa add314(s2[15], a[14]&b[3], c3[13], s3[14], c3[14]);
	fa add315(s2[16], a[15]&b[3], c3[14], s3[15], c3[15]);
	fa add316(s2[17], a[16]&b[3], c3[15], s3[16], c3[16]);
	fa add317(s2[18], a[17]&b[3], c3[16], s3[17], c3[17]);
	fa add318(s2[19], a[18]&b[3], c3[17], s3[18], c3[18]);
	fa add319(s2[20], a[19]&b[3], c3[18], s3[19], c3[19]);
	fa add320(s2[21], a[20]&b[3], c3[19], s3[20], c3[20]);
	fa add321(s2[22], a[21]&b[3], c3[20], s3[21], c3[21]);
	fa add322(s2[23], a[22]&b[3], c3[21], s3[22], c3[22]);
	fa add323(s2[24], a[23]&b[3], c3[22], s3[23], c3[23]);
	fa add324(s2[25], a[24]&b[3], c3[23], s3[24], c3[24]);
	fa add325(s2[26], a[25]&b[3], c3[24], s3[25], c3[25]);
	fa add326(s2[27], a[26]&b[3], c3[25], s3[26], c3[26]);
	fa add327(s2[28], a[27]&b[3], c3[26], s3[27], c3[27]);
	fa add328(s2[29], a[28]&b[3], c3[27], s3[28], c3[28]);
	fa add329(s2[30], a[29]&b[3], c3[28], s3[29], c3[29]);
	fa add330(s2[31], a[30]&b[3], c3[29], s3[30], c3[30]);
	fa add331(0, a[31]&b[3], c3[30], s3[31], c3[31]);
	
	
	wire [width-1:0] c4, s4;

	fa add400(s3[1], a[0]&b[4], 0, prod[4], c4[0]);
	fa add401(s3[2], a[1]&b[4], c4[0], s4[1], c4[1]);
	fa add402(s3[3], a[2]&b[4], c4[1], s4[2], c4[2]);
	fa add403(s3[4], a[3]&b[4], c4[2], s4[3], c4[3]);
	fa add404(s3[5], a[4]&b[4], c4[3], s4[4], c4[4]);
	fa add405(s3[6], a[5]&b[4], c4[4], s4[5], c4[5]);
	fa add406(s3[7], a[6]&b[4], c4[5], s4[6], c4[6]);
	fa add407(s3[8], a[7]&b[4], c4[6], s4[7], c4[7]);
	fa add408(s3[9], a[8]&b[4], c4[7], s4[8], c4[8]);
	fa add409(s3[10], a[9]&b[4], c4[8], s4[9], c4[9]);
	fa add410(s3[11], a[10]&b[4], c4[9], s4[10], c4[10]);
	fa add411(s3[12], a[11]&b[4], c4[10], s4[11], c4[11]);
	fa add412(s3[13], a[12]&b[4], c4[11], s4[12], c4[12]);
	fa add413(s3[14], a[13]&b[4], c4[12], s4[13], c4[13]);
	fa add414(s3[15], a[14]&b[4], c4[13], s4[14], c4[14]);
	fa add415(s3[16], a[15]&b[4], c4[14], s4[15], c4[15]);
	fa add416(s3[17], a[16]&b[4], c4[15], s4[16], c4[16]);
	fa add417(s3[18], a[17]&b[4], c4[16], s4[17], c4[17]);
	fa add418(s3[19], a[18]&b[4], c4[17], s4[18], c4[18]);
	fa add419(s3[20], a[19]&b[4], c4[18], s4[19], c4[19]);
	fa add420(s3[21], a[20]&b[4], c4[19], s4[20], c4[20]);
	fa add421(s3[22], a[21]&b[4], c4[20], s4[21], c4[21]);
	fa add422(s3[23], a[22]&b[4], c4[21], s4[22], c4[22]);
	fa add423(s3[24], a[23]&b[4], c4[22], s4[23], c4[23]);
	fa add424(s3[25], a[24]&b[4], c4[23], s4[24], c4[24]);
	fa add425(s3[26], a[25]&b[4], c4[24], s4[25], c4[25]);
	fa add426(s3[27], a[26]&b[4], c4[25], s4[26], c4[26]);
	fa add427(s3[28], a[27]&b[4], c4[26], s4[27], c4[27]);
	fa add428(s3[29], a[28]&b[4], c4[27], s4[28], c4[28]);
	fa add429(s3[30], a[29]&b[4], c4[28], s4[29], c4[29]);
	fa add430(s3[31], a[30]&b[4], c4[29], s4[30], c4[30]);
	fa add431(0, a[31]&b[4], c4[30], s4[31], c4[31]);
	
	
	wire [width-1:0] c5, s5;

	fa add500(s4[1], a[0]&b[5], 0, prod[5], c5[0]);
	fa add501(s4[2], a[1]&b[5], c5[0], s5[1], c5[1]);
	fa add502(s4[3], a[2]&b[5], c5[1], s5[2], c5[2]);
	fa add503(s4[4], a[3]&b[5], c5[2], s5[3], c5[3]);
	fa add504(s4[5], a[4]&b[5], c5[3], s5[4], c5[4]);
	fa add505(s4[6], a[5]&b[5], c5[4], s5[5], c5[5]);
	fa add506(s4[7], a[6]&b[5], c5[5], s5[6], c5[6]);
	fa add507(s4[8], a[7]&b[5], c5[6], s5[7], c5[7]);
	fa add508(s4[9], a[8]&b[5], c5[7], s5[8], c5[8]);
	fa add509(s4[10], a[9]&b[5], c5[8], s5[9], c5[9]);
	fa add510(s4[11], a[10]&b[5], c5[9], s5[10], c5[10]);
	fa add511(s4[12], a[11]&b[5], c5[10], s5[11], c5[11]);
	fa add512(s4[13], a[12]&b[5], c5[11], s5[12], c5[12]);
	fa add513(s4[14], a[13]&b[5], c5[12], s5[13], c5[13]);
	fa add514(s4[15], a[14]&b[5], c5[13], s5[14], c5[14]);
	fa add515(s4[16], a[15]&b[5], c5[14], s5[15], c5[15]);
	fa add516(s4[17], a[16]&b[5], c5[15], s5[16], c5[16]);
	fa add517(s4[18], a[17]&b[5], c5[16], s5[17], c5[17]);
	fa add518(s4[19], a[18]&b[5], c5[17], s5[18], c5[18]);
	fa add519(s4[20], a[19]&b[5], c5[18], s5[19], c5[19]);
	fa add520(s4[21], a[20]&b[5], c5[19], s5[20], c5[20]);
	fa add521(s4[22], a[21]&b[5], c5[20], s5[21], c5[21]);
	fa add522(s4[23], a[22]&b[5], c5[21], s5[22], c5[22]);
	fa add523(s4[24], a[23]&b[5], c5[22], s5[23], c5[23]);
	fa add524(s4[25], a[24]&b[5], c5[23], s5[24], c5[24]);
	fa add525(s4[26], a[25]&b[5], c5[24], s5[25], c5[25]);
	fa add526(s4[27], a[26]&b[5], c5[25], s5[26], c5[26]);
	fa add527(s4[28], a[27]&b[5], c5[26], s5[27], c5[27]);
	fa add528(s4[29], a[28]&b[5], c5[27], s5[28], c5[28]);
	fa add529(s4[30], a[29]&b[5], c5[28], s5[29], c5[29]);
	fa add530(s4[31], a[30]&b[5], c5[29], s5[30], c5[30]);
	fa add531(0, a[31]&b[5], c5[30], s5[31], c5[31]);
	
	
	wire [width-1:0] c6, s6;

	fa add600(s5[1], a[0]&b[6], 0, prod[6], c6[0]);
	fa add601(s5[2], a[1]&b[6], c6[0], s6[1], c6[1]);
	fa add602(s5[3], a[2]&b[6], c6[1], s6[2], c6[2]);
	fa add603(s5[4], a[3]&b[6], c6[2], s6[3], c6[3]);
	fa add604(s5[5], a[4]&b[6], c6[3], s6[4], c6[4]);
	fa add605(s5[6], a[5]&b[6], c6[4], s6[5], c6[5]);
	fa add606(s5[7], a[6]&b[6], c6[5], s6[6], c6[6]);
	fa add607(s5[8], a[7]&b[6], c6[6], s6[7], c6[7]);
	fa add608(s5[9], a[8]&b[6], c6[7], s6[8], c6[8]);
	fa add609(s5[10], a[9]&b[6], c6[8], s6[9], c6[9]);
	fa add610(s5[11], a[10]&b[6], c6[9], s6[10], c6[10]);
	fa add611(s5[12], a[11]&b[6], c6[10], s6[11], c6[11]);
	fa add612(s5[13], a[12]&b[6], c6[11], s6[12], c6[12]);
	fa add613(s5[14], a[13]&b[6], c6[12], s6[13], c6[13]);
	fa add614(s5[15], a[14]&b[6], c6[13], s6[14], c6[14]);
	fa add615(s5[16], a[15]&b[6], c6[14], s6[15], c6[15]);
	fa add616(s5[17], a[16]&b[6], c6[15], s6[16], c6[16]);
	fa add617(s5[18], a[17]&b[6], c6[16], s6[17], c6[17]);
	fa add618(s5[19], a[18]&b[6], c6[17], s6[18], c6[18]);
	fa add619(s5[20], a[19]&b[6], c6[18], s6[19], c6[19]);
	fa add620(s5[21], a[20]&b[6], c6[19], s6[20], c6[20]);
	fa add621(s5[22], a[21]&b[6], c6[20], s6[21], c6[21]);
	fa add622(s5[23], a[22]&b[6], c6[21], s6[22], c6[22]);
	fa add623(s5[24], a[23]&b[6], c6[22], s6[23], c6[23]);
	fa add624(s5[25], a[24]&b[6], c6[23], s6[24], c6[24]);
	fa add625(s5[26], a[25]&b[6], c6[24], s6[25], c6[25]);
	fa add626(s5[27], a[26]&b[6], c6[25], s6[26], c6[26]);
	fa add627(s5[28], a[27]&b[6], c6[26], s6[27], c6[27]);
	fa add628(s5[29], a[28]&b[6], c6[27], s6[28], c6[28]);
	fa add629(s5[30], a[29]&b[6], c6[28], s6[29], c6[29]);
	fa add630(s5[31], a[30]&b[6], c6[29], s6[30], c6[30]);
	fa add631(0, a[31]&b[6], c6[30], s6[31], c6[31]);
	
	
	wire [width-1:0] c7, s7;

	fa add700(s6[1], a[0]&b[7], 0, prod[7], c7[0]);
	fa add701(s6[2], a[1]&b[7], c7[0], s7[1], c7[1]);
	fa add702(s6[3], a[2]&b[7], c7[1], s7[2], c7[2]);
	fa add703(s6[4], a[3]&b[7], c7[2], s7[3], c7[3]);
	fa add704(s6[5], a[4]&b[7], c7[3], s7[4], c7[4]);
	fa add705(s6[6], a[5]&b[7], c7[4], s7[5], c7[5]);
	fa add706(s6[7], a[6]&b[7], c7[5], s7[6], c7[6]);
	fa add707(s6[8], a[7]&b[7], c7[6], s7[7], c7[7]);
	fa add708(s6[9], a[8]&b[7], c7[7], s7[8], c7[8]);
	fa add709(s6[10], a[9]&b[7], c7[8], s7[9], c7[9]);
	fa add710(s6[11], a[10]&b[7], c7[9], s7[10], c7[10]);
	fa add711(s6[12], a[11]&b[7], c7[10], s7[11], c7[11]);
	fa add712(s6[13], a[12]&b[7], c7[11], s7[12], c7[12]);
	fa add713(s6[14], a[13]&b[7], c7[12], s7[13], c7[13]);
	fa add714(s6[15], a[14]&b[7], c7[13], s7[14], c7[14]);
	fa add715(s6[16], a[15]&b[7], c7[14], s7[15], c7[15]);
	fa add716(s6[17], a[16]&b[7], c7[15], s7[16], c7[16]);
	fa add717(s6[18], a[17]&b[7], c7[16], s7[17], c7[17]);
	fa add718(s6[19], a[18]&b[7], c7[17], s7[18], c7[18]);
	fa add719(s6[20], a[19]&b[7], c7[18], s7[19], c7[19]);
	fa add720(s6[21], a[20]&b[7], c7[19], s7[20], c7[20]);
	fa add721(s6[22], a[21]&b[7], c7[20], s7[21], c7[21]);
	fa add722(s6[23], a[22]&b[7], c7[21], s7[22], c7[22]);
	fa add723(s6[24], a[23]&b[7], c7[22], s7[23], c7[23]);
	fa add724(s6[25], a[24]&b[7], c7[23], s7[24], c7[24]);
	fa add725(s6[26], a[25]&b[7], c7[24], s7[25], c7[25]);
	fa add726(s6[27], a[26]&b[7], c7[25], s7[26], c7[26]);
	fa add727(s6[28], a[27]&b[7], c7[26], s7[27], c7[27]);
	fa add728(s6[29], a[28]&b[7], c7[27], s7[28], c7[28]);
	fa add729(s6[30], a[29]&b[7], c7[28], s7[29], c7[29]);
	fa add730(s6[31], a[30]&b[7], c7[29], s7[30], c7[30]);
	fa add731(0, a[31]&b[7], c7[30], s7[31], c7[31]);
	
	
	wire [width-1:0] c8, s8;

	fa add800(s7[1], a[0]&b[8], 0, prod[8], c8[0]);
	fa add801(s7[2], a[1]&b[8], c8[0], s8[1], c8[1]);
	fa add802(s7[3], a[2]&b[8], c8[1], s8[2], c8[2]);
	fa add803(s7[4], a[3]&b[8], c8[2], s8[3], c8[3]);
	fa add804(s7[5], a[4]&b[8], c8[3], s8[4], c8[4]);
	fa add805(s7[6], a[5]&b[8], c8[4], s8[5], c8[5]);
	fa add806(s7[7], a[6]&b[8], c8[5], s8[6], c8[6]);
	fa add807(s7[8], a[7]&b[8], c8[6], s8[7], c8[7]);
	fa add808(s7[9], a[8]&b[8], c8[7], s8[8], c8[8]);
	fa add809(s7[10], a[9]&b[8], c8[8], s8[9], c8[9]);
	fa add810(s7[11], a[10]&b[8], c8[9], s8[10], c8[10]);
	fa add811(s7[12], a[11]&b[8], c8[10], s8[11], c8[11]);
	fa add812(s7[13], a[12]&b[8], c8[11], s8[12], c8[12]);
	fa add813(s7[14], a[13]&b[8], c8[12], s8[13], c8[13]);
	fa add814(s7[15], a[14]&b[8], c8[13], s8[14], c8[14]);
	fa add815(s7[16], a[15]&b[8], c8[14], s8[15], c8[15]);
	fa add816(s7[17], a[16]&b[8], c8[15], s8[16], c8[16]);
	fa add817(s7[18], a[17]&b[8], c8[16], s8[17], c8[17]);
	fa add818(s7[19], a[18]&b[8], c8[17], s8[18], c8[18]);
	fa add819(s7[20], a[19]&b[8], c8[18], s8[19], c8[19]);
	fa add820(s7[21], a[20]&b[8], c8[19], s8[20], c8[20]);
	fa add821(s7[22], a[21]&b[8], c8[20], s8[21], c8[21]);
	fa add822(s7[23], a[22]&b[8], c8[21], s8[22], c8[22]);
	fa add823(s7[24], a[23]&b[8], c8[22], s8[23], c8[23]);
	fa add824(s7[25], a[24]&b[8], c8[23], s8[24], c8[24]);
	fa add825(s7[26], a[25]&b[8], c8[24], s8[25], c8[25]);
	fa add826(s7[27], a[26]&b[8], c8[25], s8[26], c8[26]);
	fa add827(s7[28], a[27]&b[8], c8[26], s8[27], c8[27]);
	fa add828(s7[29], a[28]&b[8], c8[27], s8[28], c8[28]);
	fa add829(s7[30], a[29]&b[8], c8[28], s8[29], c8[29]);
	fa add830(s7[31], a[30]&b[8], c8[29], s8[30], c8[30]);
	fa add831(0, a[31]&b[8], c8[30], s8[31], c8[31]);
	
	
	wire [width-1:0] c9, s9;

	fa add900(s8[1], a[0]&b[9], 0, prod[9], c9[0]);
	fa add901(s8[2], a[1]&b[9], c9[0], s9[1], c9[1]);
	fa add902(s8[3], a[2]&b[9], c9[1], s9[2], c9[2]);
	fa add903(s8[4], a[3]&b[9], c9[2], s9[3], c9[3]);
	fa add904(s8[5], a[4]&b[9], c9[3], s9[4], c9[4]);
	fa add905(s8[6], a[5]&b[9], c9[4], s9[5], c9[5]);
	fa add906(s8[7], a[6]&b[9], c9[5], s9[6], c9[6]);
	fa add907(s8[8], a[7]&b[9], c9[6], s9[7], c9[7]);
	fa add908(s8[9], a[8]&b[9], c9[7], s9[8], c9[8]);
	fa add909(s8[10], a[9]&b[9], c9[8], s9[9], c9[9]);
	fa add910(s8[11], a[10]&b[9], c9[9], s9[10], c9[10]);
	fa add911(s8[12], a[11]&b[9], c9[10], s9[11], c9[11]);
	fa add912(s8[13], a[12]&b[9], c9[11], s9[12], c9[12]);
	fa add913(s8[14], a[13]&b[9], c9[12], s9[13], c9[13]);
	fa add914(s8[15], a[14]&b[9], c9[13], s9[14], c9[14]);
	fa add915(s8[16], a[15]&b[9], c9[14], s9[15], c9[15]);
	fa add916(s8[17], a[16]&b[9], c9[15], s9[16], c9[16]);
	fa add917(s8[18], a[17]&b[9], c9[16], s9[17], c9[17]);
	fa add918(s8[19], a[18]&b[9], c9[17], s9[18], c9[18]);
	fa add919(s8[20], a[19]&b[9], c9[18], s9[19], c9[19]);
	fa add920(s8[21], a[20]&b[9], c9[19], s9[20], c9[20]);
	fa add921(s8[22], a[21]&b[9], c9[20], s9[21], c9[21]);
	fa add922(s8[23], a[22]&b[9], c9[21], s9[22], c9[22]);
	fa add923(s8[24], a[23]&b[9], c9[22], s9[23], c9[23]);
	fa add924(s8[25], a[24]&b[9], c9[23], s9[24], c9[24]);
	fa add925(s8[26], a[25]&b[9], c9[24], s9[25], c9[25]);
	fa add926(s8[27], a[26]&b[9], c9[25], s9[26], c9[26]);
	fa add927(s8[28], a[27]&b[9], c9[26], s9[27], c9[27]);
	fa add928(s8[29], a[28]&b[9], c9[27], s9[28], c9[28]);
	fa add929(s8[30], a[29]&b[9], c9[28], s9[29], c9[29]);
	fa add930(s8[31], a[30]&b[9], c9[29], s9[30], c9[30]);
	fa add931(0, a[31]&b[9], c9[30], s9[31], c9[31]);
	
	
	wire [width-1:0] c10, s10;

	fa add1000(s9[1], a[0]&b[10], 0, prod[10], c10[0]);
	fa add1001(s9[2], a[1]&b[10], c10[0], s10[1], c10[1]);
	fa add1002(s9[3], a[2]&b[10], c10[1], s10[2], c10[2]);
	fa add1003(s9[4], a[3]&b[10], c10[2], s10[3], c10[3]);
	fa add1004(s9[5], a[4]&b[10], c10[3], s10[4], c10[4]);
	fa add1005(s9[6], a[5]&b[10], c10[4], s10[5], c10[5]);
	fa add1006(s9[7], a[6]&b[10], c10[5], s10[6], c10[6]);
	fa add1007(s9[8], a[7]&b[10], c10[6], s10[7], c10[7]);
	fa add1008(s9[9], a[8]&b[10], c10[7], s10[8], c10[8]);
	fa add1009(s9[10], a[9]&b[10], c10[8], s10[9], c10[9]);
	fa add1010(s9[11], a[10]&b[10], c10[9], s10[10], c10[10]);
	fa add1011(s9[12], a[11]&b[10], c10[10], s10[11], c10[11]);
	fa add1012(s9[13], a[12]&b[10], c10[11], s10[12], c10[12]);
	fa add1013(s9[14], a[13]&b[10], c10[12], s10[13], c10[13]);
	fa add1014(s9[15], a[14]&b[10], c10[13], s10[14], c10[14]);
	fa add1015(s9[16], a[15]&b[10], c10[14], s10[15], c10[15]);
	fa add1016(s9[17], a[16]&b[10], c10[15], s10[16], c10[16]);
	fa add1017(s9[18], a[17]&b[10], c10[16], s10[17], c10[17]);
	fa add1018(s9[19], a[18]&b[10], c10[17], s10[18], c10[18]);
	fa add1019(s9[20], a[19]&b[10], c10[18], s10[19], c10[19]);
	fa add1020(s9[21], a[20]&b[10], c10[19], s10[20], c10[20]);
	fa add1021(s9[22], a[21]&b[10], c10[20], s10[21], c10[21]);
	fa add1022(s9[23], a[22]&b[10], c10[21], s10[22], c10[22]);
	fa add1023(s9[24], a[23]&b[10], c10[22], s10[23], c10[23]);
	fa add1024(s9[25], a[24]&b[10], c10[23], s10[24], c10[24]);
	fa add1025(s9[26], a[25]&b[10], c10[24], s10[25], c10[25]);
	fa add1026(s9[27], a[26]&b[10], c10[25], s10[26], c10[26]);
	fa add1027(s9[28], a[27]&b[10], c10[26], s10[27], c10[27]);
	fa add1028(s9[29], a[28]&b[10], c10[27], s10[28], c10[28]);
	fa add1029(s9[30], a[29]&b[10], c10[28], s10[29], c10[29]);
	fa add1030(s9[31], a[30]&b[10], c10[29], s10[30], c10[30]);
	fa add1031(0, a[31]&b[10], c10[30], s10[31], c10[31]);
		
	
	wire [width-1:0] c11, s11;

	fa add1100(s10[1], a[0]&b[11], 0, prod[11], c11[0]);
	fa add1101(s10[2], a[1]&b[11], c11[0], s11[1], c11[1]);
	fa add1102(s10[3], a[2]&b[11], c11[1], s11[2], c11[2]);
	fa add1103(s10[4], a[3]&b[11], c11[2], s11[3], c11[3]);
	fa add1104(s10[5], a[4]&b[11], c11[3], s11[4], c11[4]);
	fa add1105(s10[6], a[5]&b[11], c11[4], s11[5], c11[5]);
	fa add1106(s10[7], a[6]&b[11], c11[5], s11[6], c11[6]);
	fa add1107(s10[8], a[7]&b[11], c11[6], s11[7], c11[7]);
	fa add1108(s10[9], a[8]&b[11], c11[7], s11[8], c11[8]);
	fa add1109(s10[10], a[9]&b[11], c11[8], s11[9], c11[9]);
	fa add1110(s10[11], a[10]&b[11], c11[9], s11[10], c11[10]);
	fa add1111(s10[12], a[11]&b[11], c11[10], s11[11], c11[11]);
	fa add1112(s10[13], a[12]&b[11], c11[11], s11[12], c11[12]);
	fa add1113(s10[14], a[13]&b[11], c11[12], s11[13], c11[13]);
	fa add1114(s10[15], a[14]&b[11], c11[13], s11[14], c11[14]);
	fa add1115(s10[16], a[15]&b[11], c11[14], s11[15], c11[15]);
	fa add1116(s10[17], a[16]&b[11], c11[15], s11[16], c11[16]);
	fa add1117(s10[18], a[17]&b[11], c11[16], s11[17], c11[17]);
	fa add1118(s10[19], a[18]&b[11], c11[17], s11[18], c11[18]);
	fa add1119(s10[20], a[19]&b[11], c11[18], s11[19], c11[19]);
	fa add1120(s10[21], a[20]&b[11], c11[19], s11[20], c11[20]);
	fa add1121(s10[22], a[21]&b[11], c11[20], s11[21], c11[21]);
	fa add1122(s10[23], a[22]&b[11], c11[21], s11[22], c11[22]);
	fa add1123(s10[24], a[23]&b[11], c11[22], s11[23], c11[23]);
	fa add1124(s10[25], a[24]&b[11], c11[23], s11[24], c11[24]);
	fa add1125(s10[26], a[25]&b[11], c11[24], s11[25], c11[25]);
	fa add1126(s10[27], a[26]&b[11], c11[25], s11[26], c11[26]);
	fa add1127(s10[28], a[27]&b[11], c11[26], s11[27], c11[27]);
	fa add1128(s10[29], a[28]&b[11], c11[27], s11[28], c11[28]);
	fa add1129(s10[30], a[29]&b[11], c11[28], s11[29], c11[29]);
	fa add1130(s10[31], a[30]&b[11], c11[29], s11[30], c11[30]);
	fa add1131(0, a[31]&b[11], c11[30], s11[31], c11[31]);
		
	
	wire [width-1:0] c12, s12;

	fa add1200(s11[1], a[0]&b[12], 0, prod[12], c12[0]);
	fa add1201(s11[2], a[1]&b[12], c12[0], s12[1], c12[1]);
	fa add1202(s11[3], a[2]&b[12], c12[1], s12[2], c12[2]);
	fa add1203(s11[4], a[3]&b[12], c12[2], s12[3], c12[3]);
	fa add1204(s11[5], a[4]&b[12], c12[3], s12[4], c12[4]);
	fa add1205(s11[6], a[5]&b[12], c12[4], s12[5], c12[5]);
	fa add1206(s11[7], a[6]&b[12], c12[5], s12[6], c12[6]);
	fa add1207(s11[8], a[7]&b[12], c12[6], s12[7], c12[7]);
	fa add1208(s11[9], a[8]&b[12], c12[7], s12[8], c12[8]);
	fa add1209(s11[10], a[9]&b[12], c12[8], s12[9], c12[9]);
	fa add1210(s11[11], a[10]&b[12], c12[9], s12[10], c12[10]);
	fa add1211(s11[12], a[11]&b[12], c12[10], s12[11], c12[11]);
	fa add1212(s11[13], a[12]&b[12], c12[11], s12[12], c12[12]);
	fa add1213(s11[14], a[13]&b[12], c12[12], s12[13], c12[13]);
	fa add1214(s11[15], a[14]&b[12], c12[13], s12[14], c12[14]);
	fa add1215(s11[16], a[15]&b[12], c12[14], s12[15], c12[15]);
	fa add1216(s11[17], a[16]&b[12], c12[15], s12[16], c12[16]);
	fa add1217(s11[18], a[17]&b[12], c12[16], s12[17], c12[17]);
	fa add1218(s11[19], a[18]&b[12], c12[17], s12[18], c12[18]);
	fa add1219(s11[20], a[19]&b[12], c12[18], s12[19], c12[19]);
	fa add1220(s11[21], a[20]&b[12], c12[19], s12[20], c12[20]);
	fa add1221(s11[22], a[21]&b[12], c12[20], s12[21], c12[21]);
	fa add1222(s11[23], a[22]&b[12], c12[21], s12[22], c12[22]);
	fa add1223(s11[24], a[23]&b[12], c12[22], s12[23], c12[23]);
	fa add1224(s11[25], a[24]&b[12], c12[23], s12[24], c12[24]);
	fa add1225(s11[26], a[25]&b[12], c12[24], s12[25], c12[25]);
	fa add1226(s11[27], a[26]&b[12], c12[25], s12[26], c12[26]);
	fa add1227(s11[28], a[27]&b[12], c12[26], s12[27], c12[27]);
	fa add1228(s11[29], a[28]&b[12], c12[27], s12[28], c12[28]);
	fa add1229(s11[30], a[29]&b[12], c12[28], s12[29], c12[29]);
	fa add1230(s11[31], a[30]&b[12], c12[29], s12[30], c12[30]);
	fa add1231(0, a[31]&b[12], c12[30], s12[31], c12[31]);
		
	
	wire [width-1:0] c13, s13;

	fa add1300(s12[1], a[0]&b[13], 0, prod[13], c13[0]);
	fa add1301(s12[2], a[1]&b[13], c13[0], s13[1], c13[1]);
	fa add1302(s12[3], a[2]&b[13], c13[1], s13[2], c13[2]);
	fa add1303(s12[4], a[3]&b[13], c13[2], s13[3], c13[3]);
	fa add1304(s12[5], a[4]&b[13], c13[3], s13[4], c13[4]);
	fa add1305(s12[6], a[5]&b[13], c13[4], s13[5], c13[5]);
	fa add1306(s12[7], a[6]&b[13], c13[5], s13[6], c13[6]);
	fa add1307(s12[8], a[7]&b[13], c13[6], s13[7], c13[7]);
	fa add1308(s12[9], a[8]&b[13], c13[7], s13[8], c13[8]);
	fa add1309(s12[10], a[9]&b[13], c13[8], s13[9], c13[9]);
	fa add1310(s12[11], a[10]&b[13], c13[9], s13[10], c13[10]);
	fa add1311(s12[12], a[11]&b[13], c13[10], s13[11], c13[11]);
	fa add1312(s12[13], a[12]&b[13], c13[11], s13[12], c13[12]);
	fa add1313(s12[14], a[13]&b[13], c13[12], s13[13], c13[13]);
	fa add1314(s12[15], a[14]&b[13], c13[13], s13[14], c13[14]);
	fa add1315(s12[16], a[15]&b[13], c13[14], s13[15], c13[15]);
	fa add1316(s12[17], a[16]&b[13], c13[15], s13[16], c13[16]);
	fa add1317(s12[18], a[17]&b[13], c13[16], s13[17], c13[17]);
	fa add1318(s12[19], a[18]&b[13], c13[17], s13[18], c13[18]);
	fa add1319(s12[20], a[19]&b[13], c13[18], s13[19], c13[19]);
	fa add1320(s12[21], a[20]&b[13], c13[19], s13[20], c13[20]);
	fa add1321(s12[22], a[21]&b[13], c13[20], s13[21], c13[21]);
	fa add1322(s12[23], a[22]&b[13], c13[21], s13[22], c13[22]);
	fa add1323(s12[24], a[23]&b[13], c13[22], s13[23], c13[23]);
	fa add1324(s12[25], a[24]&b[13], c13[23], s13[24], c13[24]);
	fa add1325(s12[26], a[25]&b[13], c13[24], s13[25], c13[25]);
	fa add1326(s12[27], a[26]&b[13], c13[25], s13[26], c13[26]);
	fa add1327(s12[28], a[27]&b[13], c13[26], s13[27], c13[27]);
	fa add1328(s12[29], a[28]&b[13], c13[27], s13[28], c13[28]);
	fa add1329(s12[30], a[29]&b[13], c13[28], s13[29], c13[29]);
	fa add1330(s12[31], a[30]&b[13], c13[29], s13[30], c13[30]);
	fa add1331(0, a[31]&b[13], c13[30], s13[31], c13[31]);
		
	
	wire [width-1:0] c14, s14;

	fa add1400(s13[1], a[0]&b[14], 0, prod[14], c14[0]);
	fa add1401(s13[2], a[1]&b[14], c14[0], s14[1], c14[1]);
	fa add1402(s13[3], a[2]&b[14], c14[1], s14[2], c14[2]);
	fa add1403(s13[4], a[3]&b[14], c14[2], s14[3], c14[3]);
	fa add1404(s13[5], a[4]&b[14], c14[3], s14[4], c14[4]);
	fa add1405(s13[6], a[5]&b[14], c14[4], s14[5], c14[5]);
	fa add1406(s13[7], a[6]&b[14], c14[5], s14[6], c14[6]);
	fa add1407(s13[8], a[7]&b[14], c14[6], s14[7], c14[7]);
	fa add1408(s13[9], a[8]&b[14], c14[7], s14[8], c14[8]);
	fa add1409(s13[10], a[9]&b[14], c14[8], s14[9], c14[9]);
	fa add1410(s13[11], a[10]&b[14], c14[9], s14[10], c14[10]);
	fa add1411(s13[12], a[11]&b[14], c14[10], s14[11], c14[11]);
	fa add1412(s13[13], a[12]&b[14], c14[11], s14[12], c14[12]);
	fa add1413(s13[14], a[13]&b[14], c14[12], s14[13], c14[13]);
	fa add1414(s13[15], a[14]&b[14], c14[13], s14[14], c14[14]);
	fa add1415(s13[16], a[15]&b[14], c14[14], s14[15], c14[15]);
	fa add1416(s13[17], a[16]&b[14], c14[15], s14[16], c14[16]);
	fa add1417(s13[18], a[17]&b[14], c14[16], s14[17], c14[17]);
	fa add1418(s13[19], a[18]&b[14], c14[17], s14[18], c14[18]);
	fa add1419(s13[20], a[19]&b[14], c14[18], s14[19], c14[19]);
	fa add1420(s13[21], a[20]&b[14], c14[19], s14[20], c14[20]);
	fa add1421(s13[22], a[21]&b[14], c14[20], s14[21], c14[21]);
	fa add1422(s13[23], a[22]&b[14], c14[21], s14[22], c14[22]);
	fa add1423(s13[24], a[23]&b[14], c14[22], s14[23], c14[23]);
	fa add1424(s13[25], a[24]&b[14], c14[23], s14[24], c14[24]);
	fa add1425(s13[26], a[25]&b[14], c14[24], s14[25], c14[25]);
	fa add1426(s13[27], a[26]&b[14], c14[25], s14[26], c14[26]);
	fa add1427(s13[28], a[27]&b[14], c14[26], s14[27], c14[27]);
	fa add1428(s13[29], a[28]&b[14], c14[27], s14[28], c14[28]);
	fa add1429(s13[30], a[29]&b[14], c14[28], s14[29], c14[29]);
	fa add1430(s13[31], a[30]&b[14], c14[29], s14[30], c14[30]);
	fa add1431(0, a[31]&b[14], c14[30], s14[31], c14[31]);
		
	
	wire [width-1:0] c15, s15;

	fa add1500(s14[1], a[0]&b[15], 0, prod[15], c15[0]);
	fa add1501(s14[2], a[1]&b[15], c15[0], s15[1], c15[1]);
	fa add1502(s14[3], a[2]&b[15], c15[1], s15[2], c15[2]);
	fa add1503(s14[4], a[3]&b[15], c15[2], s15[3], c15[3]);
	fa add1504(s14[5], a[4]&b[15], c15[3], s15[4], c15[4]);
	fa add1505(s14[6], a[5]&b[15], c15[4], s15[5], c15[5]);
	fa add1506(s14[7], a[6]&b[15], c15[5], s15[6], c15[6]);
	fa add1507(s14[8], a[7]&b[15], c15[6], s15[7], c15[7]);
	fa add1508(s14[9], a[8]&b[15], c15[7], s15[8], c15[8]);
	fa add1509(s14[10], a[9]&b[15], c15[8], s15[9], c15[9]);
	fa add1510(s14[11], a[10]&b[15], c15[9], s15[10], c15[10]);
	fa add1511(s14[12], a[11]&b[15], c15[10], s15[11], c15[11]);
	fa add1512(s14[13], a[12]&b[15], c15[11], s15[12], c15[12]);
	fa add1513(s14[14], a[13]&b[15], c15[12], s15[13], c15[13]);
	fa add1514(s14[15], a[14]&b[15], c15[13], s15[14], c15[14]);
	fa add1515(s14[16], a[15]&b[15], c15[14], s15[15], c15[15]);
	fa add1516(s14[17], a[16]&b[15], c15[15], s15[16], c15[16]);
	fa add1517(s14[18], a[17]&b[15], c15[16], s15[17], c15[17]);
	fa add1518(s14[19], a[18]&b[15], c15[17], s15[18], c15[18]);
	fa add1519(s14[20], a[19]&b[15], c15[18], s15[19], c15[19]);
	fa add1520(s14[21], a[20]&b[15], c15[19], s15[20], c15[20]);
	fa add1521(s14[22], a[21]&b[15], c15[20], s15[21], c15[21]);
	fa add1522(s14[23], a[22]&b[15], c15[21], s15[22], c15[22]);
	fa add1523(s14[24], a[23]&b[15], c15[22], s15[23], c15[23]);
	fa add1524(s14[25], a[24]&b[15], c15[23], s15[24], c15[24]);
	fa add1525(s14[26], a[25]&b[15], c15[24], s15[25], c15[25]);
	fa add1526(s14[27], a[26]&b[15], c15[25], s15[26], c15[26]);
	fa add1527(s14[28], a[27]&b[15], c15[26], s15[27], c15[27]);
	fa add1528(s14[29], a[28]&b[15], c15[27], s15[28], c15[28]);
	fa add1529(s14[30], a[29]&b[15], c15[28], s15[29], c15[29]);
	fa add1530(s14[31], a[30]&b[15], c15[29], s15[30], c15[30]);
	fa add1531(0, a[31]&b[15], c15[30], s15[31], c15[31]);
		
	
	wire [width-1:0] c16, s16;

	fa add1600(s15[1], a[0]&b[16], 0, prod[16], c16[0]);
	fa add1601(s15[2], a[1]&b[16], c16[0], s16[1], c16[1]);
	fa add1602(s15[3], a[2]&b[16], c16[1], s16[2], c16[2]);
	fa add1603(s15[4], a[3]&b[16], c16[2], s16[3], c16[3]);
	fa add1604(s15[5], a[4]&b[16], c16[3], s16[4], c16[4]);
	fa add1605(s15[6], a[5]&b[16], c16[4], s16[5], c16[5]);
	fa add1606(s15[7], a[6]&b[16], c16[5], s16[6], c16[6]);
	fa add1607(s15[8], a[7]&b[16], c16[6], s16[7], c16[7]);
	fa add1608(s15[9], a[8]&b[16], c16[7], s16[8], c16[8]);
	fa add1609(s15[10], a[9]&b[16], c16[8], s16[9], c16[9]);
	fa add1610(s15[11], a[10]&b[16], c16[9], s16[10], c16[10]);
	fa add1611(s15[12], a[11]&b[16], c16[10], s16[11], c16[11]);
	fa add1612(s15[13], a[12]&b[16], c16[11], s16[12], c16[12]);
	fa add1613(s15[14], a[13]&b[16], c16[12], s16[13], c16[13]);
	fa add1614(s15[15], a[14]&b[16], c16[13], s16[14], c16[14]);
	fa add1615(s15[16], a[15]&b[16], c16[14], s16[15], c16[15]);
	fa add1616(s15[17], a[16]&b[16], c16[15], s16[16], c16[16]);
	fa add1617(s15[18], a[17]&b[16], c16[16], s16[17], c16[17]);
	fa add1618(s15[19], a[18]&b[16], c16[17], s16[18], c16[18]);
	fa add1619(s15[20], a[19]&b[16], c16[18], s16[19], c16[19]);
	fa add1620(s15[21], a[20]&b[16], c16[19], s16[20], c16[20]);
	fa add1621(s15[22], a[21]&b[16], c16[20], s16[21], c16[21]);
	fa add1622(s15[23], a[22]&b[16], c16[21], s16[22], c16[22]);
	fa add1623(s15[24], a[23]&b[16], c16[22], s16[23], c16[23]);
	fa add1624(s15[25], a[24]&b[16], c16[23], s16[24], c16[24]);
	fa add1625(s15[26], a[25]&b[16], c16[24], s16[25], c16[25]);
	fa add1626(s15[27], a[26]&b[16], c16[25], s16[26], c16[26]);
	fa add1627(s15[28], a[27]&b[16], c16[26], s16[27], c16[27]);
	fa add1628(s15[29], a[28]&b[16], c16[27], s16[28], c16[28]);
	fa add1629(s15[30], a[29]&b[16], c16[28], s16[29], c16[29]);
	fa add1630(s15[31], a[30]&b[16], c16[29], s16[30], c16[30]);
	fa add1631(0, a[31]&b[16], c16[30], s16[31], c16[31]);
		
	
	wire [width-1:0] c17, s17;

	fa add1700(s16[1], a[0]&b[17], 0, prod[17], c17[0]);
	fa add1701(s16[2], a[1]&b[17], c17[0], s17[1], c17[1]);
	fa add1702(s16[3], a[2]&b[17], c17[1], s17[2], c17[2]);
	fa add1703(s16[4], a[3]&b[17], c17[2], s17[3], c17[3]);
	fa add1704(s16[5], a[4]&b[17], c17[3], s17[4], c17[4]);
	fa add1705(s16[6], a[5]&b[17], c17[4], s17[5], c17[5]);
	fa add1706(s16[7], a[6]&b[17], c17[5], s17[6], c17[6]);
	fa add1707(s16[8], a[7]&b[17], c17[6], s17[7], c17[7]);
	fa add1708(s16[9], a[8]&b[17], c17[7], s17[8], c17[8]);
	fa add1709(s16[10], a[9]&b[17], c17[8], s17[9], c17[9]);
	fa add1710(s16[11], a[10]&b[17], c17[9], s17[10], c17[10]);
	fa add1711(s16[12], a[11]&b[17], c17[10], s17[11], c17[11]);
	fa add1712(s16[13], a[12]&b[17], c17[11], s17[12], c17[12]);
	fa add1713(s16[14], a[13]&b[17], c17[12], s17[13], c17[13]);
	fa add1714(s16[15], a[14]&b[17], c17[13], s17[14], c17[14]);
	fa add1715(s16[16], a[15]&b[17], c17[14], s17[15], c17[15]);
	fa add1716(s16[17], a[16]&b[17], c17[15], s17[16], c17[16]);
	fa add1717(s16[18], a[17]&b[17], c17[16], s17[17], c17[17]);
	fa add1718(s16[19], a[18]&b[17], c17[17], s17[18], c17[18]);
	fa add1719(s16[20], a[19]&b[17], c17[18], s17[19], c17[19]);
	fa add1720(s16[21], a[20]&b[17], c17[19], s17[20], c17[20]);
	fa add1721(s16[22], a[21]&b[17], c17[20], s17[21], c17[21]);
	fa add1722(s16[23], a[22]&b[17], c17[21], s17[22], c17[22]);
	fa add1723(s16[24], a[23]&b[17], c17[22], s17[23], c17[23]);
	fa add1724(s16[25], a[24]&b[17], c17[23], s17[24], c17[24]);
	fa add1725(s16[26], a[25]&b[17], c17[24], s17[25], c17[25]);
	fa add1726(s16[27], a[26]&b[17], c17[25], s17[26], c17[26]);
	fa add1727(s16[28], a[27]&b[17], c17[26], s17[27], c17[27]);
	fa add1728(s16[29], a[28]&b[17], c17[27], s17[28], c17[28]);
	fa add1729(s16[30], a[29]&b[17], c17[28], s17[29], c17[29]);
	fa add1730(s16[31], a[30]&b[17], c17[29], s17[30], c17[30]);
	fa add1731(0, a[31]&b[17], c17[30], s17[31], c17[31]);
		
	
	wire [width-1:0] c18, s18;

	fa add1800(s17[1], a[0]&b[18], 0, prod[18], c18[0]);
	fa add1801(s17[2], a[1]&b[18], c18[0], s18[1], c18[1]);
	fa add1802(s17[3], a[2]&b[18], c18[1], s18[2], c18[2]);
	fa add1803(s17[4], a[3]&b[18], c18[2], s18[3], c18[3]);
	fa add1804(s17[5], a[4]&b[18], c18[3], s18[4], c18[4]);
	fa add1805(s17[6], a[5]&b[18], c18[4], s18[5], c18[5]);
	fa add1806(s17[7], a[6]&b[18], c18[5], s18[6], c18[6]);
	fa add1807(s17[8], a[7]&b[18], c18[6], s18[7], c18[7]);
	fa add1808(s17[9], a[8]&b[18], c18[7], s18[8], c18[8]);
	fa add1809(s17[10], a[9]&b[18], c18[8], s18[9], c18[9]);
	fa add1810(s17[11], a[10]&b[18], c18[9], s18[10], c18[10]);
	fa add1811(s17[12], a[11]&b[18], c18[10], s18[11], c18[11]);
	fa add1812(s17[13], a[12]&b[18], c18[11], s18[12], c18[12]);
	fa add1813(s17[14], a[13]&b[18], c18[12], s18[13], c18[13]);
	fa add1814(s17[15], a[14]&b[18], c18[13], s18[14], c18[14]);
	fa add1815(s17[16], a[15]&b[18], c18[14], s18[15], c18[15]);
	fa add1816(s17[17], a[16]&b[18], c18[15], s18[16], c18[16]);
	fa add1817(s17[18], a[17]&b[18], c18[16], s18[17], c18[17]);
	fa add1818(s17[19], a[18]&b[18], c18[17], s18[18], c18[18]);
	fa add1819(s17[20], a[19]&b[18], c18[18], s18[19], c18[19]);
	fa add1820(s17[21], a[20]&b[18], c18[19], s18[20], c18[20]);
	fa add1821(s17[22], a[21]&b[18], c18[20], s18[21], c18[21]);
	fa add1822(s17[23], a[22]&b[18], c18[21], s18[22], c18[22]);
	fa add1823(s17[24], a[23]&b[18], c18[22], s18[23], c18[23]);
	fa add1824(s17[25], a[24]&b[18], c18[23], s18[24], c18[24]);
	fa add1825(s17[26], a[25]&b[18], c18[24], s18[25], c18[25]);
	fa add1826(s17[27], a[26]&b[18], c18[25], s18[26], c18[26]);
	fa add1827(s17[28], a[27]&b[18], c18[26], s18[27], c18[27]);
	fa add1828(s17[29], a[28]&b[18], c18[27], s18[28], c18[28]);
	fa add1829(s17[30], a[29]&b[18], c18[28], s18[29], c18[29]);
	fa add1830(s17[31], a[30]&b[18], c18[29], s18[30], c18[30]);
	fa add1831(0, a[31]&b[18], c18[30], s18[31], c18[31]);
		
	
	wire [width-1:0] c19, s19;

	fa add1900(s18[1], a[0]&b[19], 0, prod[19], c19[0]);
	fa add1901(s18[2], a[1]&b[19], c19[0], s19[1], c19[1]);
	fa add1902(s18[3], a[2]&b[19], c19[1], s19[2], c19[2]);
	fa add1903(s18[4], a[3]&b[19], c19[2], s19[3], c19[3]);
	fa add1904(s18[5], a[4]&b[19], c19[3], s19[4], c19[4]);
	fa add1905(s18[6], a[5]&b[19], c19[4], s19[5], c19[5]);
	fa add1906(s18[7], a[6]&b[19], c19[5], s19[6], c19[6]);
	fa add1907(s18[8], a[7]&b[19], c19[6], s19[7], c19[7]);
	fa add1908(s18[9], a[8]&b[19], c19[7], s19[8], c19[8]);
	fa add1909(s18[10], a[9]&b[19], c19[8], s19[9], c19[9]);
	fa add1910(s18[11], a[10]&b[19], c19[9], s19[10], c19[10]);
	fa add1911(s18[12], a[11]&b[19], c19[10], s19[11], c19[11]);
	fa add1912(s18[13], a[12]&b[19], c19[11], s19[12], c19[12]);
	fa add1913(s18[14], a[13]&b[19], c19[12], s19[13], c19[13]);
	fa add1914(s18[15], a[14]&b[19], c19[13], s19[14], c19[14]);
	fa add1915(s18[16], a[15]&b[19], c19[14], s19[15], c19[15]);
	fa add1916(s18[17], a[16]&b[19], c19[15], s19[16], c19[16]);
	fa add1917(s18[18], a[17]&b[19], c19[16], s19[17], c19[17]);
	fa add1918(s18[19], a[18]&b[19], c19[17], s19[18], c19[18]);
	fa add1919(s18[20], a[19]&b[19], c19[18], s19[19], c19[19]);
	fa add1920(s18[21], a[20]&b[19], c19[19], s19[20], c19[20]);
	fa add1921(s18[22], a[21]&b[19], c19[20], s19[21], c19[21]);
	fa add1922(s18[23], a[22]&b[19], c19[21], s19[22], c19[22]);
	fa add1923(s18[24], a[23]&b[19], c19[22], s19[23], c19[23]);
	fa add1924(s18[25], a[24]&b[19], c19[23], s19[24], c19[24]);
	fa add1925(s18[26], a[25]&b[19], c19[24], s19[25], c19[25]);
	fa add1926(s18[27], a[26]&b[19], c19[25], s19[26], c19[26]);
	fa add1927(s18[28], a[27]&b[19], c19[26], s19[27], c19[27]);
	fa add1928(s18[29], a[28]&b[19], c19[27], s19[28], c19[28]);
	fa add1929(s18[30], a[29]&b[19], c19[28], s19[29], c19[29]);
	fa add1930(s18[31], a[30]&b[19], c19[29], s19[30], c19[30]);
	fa add1931(0, a[31]&b[19], c19[30], s19[31], c19[31]);
		
	
	wire [width-1:0] c20, s20;

	fa add2000(s19[1], a[0]&b[20], 0, prod[20], c20[0]);
	fa add2001(s19[2], a[1]&b[20], c20[0], s20[1], c20[1]);
	fa add2002(s19[3], a[2]&b[20], c20[1], s20[2], c20[2]);
	fa add2003(s19[4], a[3]&b[20], c20[2], s20[3], c20[3]);
	fa add2004(s19[5], a[4]&b[20], c20[3], s20[4], c20[4]);
	fa add2005(s19[6], a[5]&b[20], c20[4], s20[5], c20[5]);
	fa add2006(s19[7], a[6]&b[20], c20[5], s20[6], c20[6]);
	fa add2007(s19[8], a[7]&b[20], c20[6], s20[7], c20[7]);
	fa add2008(s19[9], a[8]&b[20], c20[7], s20[8], c20[8]);
	fa add2009(s19[10], a[9]&b[20], c20[8], s20[9], c20[9]);
	fa add2010(s19[11], a[10]&b[20], c20[9], s20[10], c20[10]);
	fa add2011(s19[12], a[11]&b[20], c20[10], s20[11], c20[11]);
	fa add2012(s19[13], a[12]&b[20], c20[11], s20[12], c20[12]);
	fa add2013(s19[14], a[13]&b[20], c20[12], s20[13], c20[13]);
	fa add2014(s19[15], a[14]&b[20], c20[13], s20[14], c20[14]);
	fa add2015(s19[16], a[15]&b[20], c20[14], s20[15], c20[15]);
	fa add2016(s19[17], a[16]&b[20], c20[15], s20[16], c20[16]);
	fa add2017(s19[18], a[17]&b[20], c20[16], s20[17], c20[17]);
	fa add2018(s19[19], a[18]&b[20], c20[17], s20[18], c20[18]);
	fa add2019(s19[20], a[19]&b[20], c20[18], s20[19], c20[19]);
	fa add2020(s19[21], a[20]&b[20], c20[19], s20[20], c20[20]);
	fa add2021(s19[22], a[21]&b[20], c20[20], s20[21], c20[21]);
	fa add2022(s19[23], a[22]&b[20], c20[21], s20[22], c20[22]);
	fa add2023(s19[24], a[23]&b[20], c20[22], s20[23], c20[23]);
	fa add2024(s19[25], a[24]&b[20], c20[23], s20[24], c20[24]);
	fa add2025(s19[26], a[25]&b[20], c20[24], s20[25], c20[25]);
	fa add2026(s19[27], a[26]&b[20], c20[25], s20[26], c20[26]);
	fa add2027(s19[28], a[27]&b[20], c20[26], s20[27], c20[27]);
	fa add2028(s19[29], a[28]&b[20], c20[27], s20[28], c20[28]);
	fa add2029(s19[30], a[29]&b[20], c20[28], s20[29], c20[29]);
	fa add2030(s19[31], a[30]&b[20], c20[29], s20[30], c20[30]);
	fa add2031(0, a[31]&b[20], c20[30], s20[31], c20[31]);
	
		
	
	wire [width-1:0] c21, s21;

	fa add2100(s20[1], a[0]&b[21], 0, prod[21], c21[0]);
	fa add2101(s20[2], a[1]&b[21], c21[0], s21[1], c21[1]);
	fa add2102(s20[3], a[2]&b[21], c21[1], s21[2], c21[2]);
	fa add2103(s20[4], a[3]&b[21], c21[2], s21[3], c21[3]);
	fa add2104(s20[5], a[4]&b[21], c21[3], s21[4], c21[4]);
	fa add2105(s20[6], a[5]&b[21], c21[4], s21[5], c21[5]);
	fa add2106(s20[7], a[6]&b[21], c21[5], s21[6], c21[6]);
	fa add2107(s20[8], a[7]&b[21], c21[6], s21[7], c21[7]);
	fa add2108(s20[9], a[8]&b[21], c21[7], s21[8], c21[8]);
	fa add2109(s20[10], a[9]&b[21], c21[8], s21[9], c21[9]);
	fa add2110(s20[11], a[10]&b[21], c21[9], s21[10], c21[10]);
	fa add2111(s20[12], a[11]&b[21], c21[10], s21[11], c21[11]);
	fa add2112(s20[13], a[12]&b[21], c21[11], s21[12], c21[12]);
	fa add2113(s20[14], a[13]&b[21], c21[12], s21[13], c21[13]);
	fa add2114(s20[15], a[14]&b[21], c21[13], s21[14], c21[14]);
	fa add2115(s20[16], a[15]&b[21], c21[14], s21[15], c21[15]);
	fa add2116(s20[17], a[16]&b[21], c21[15], s21[16], c21[16]);
	fa add2117(s20[18], a[17]&b[21], c21[16], s21[17], c21[17]);
	fa add2118(s20[19], a[18]&b[21], c21[17], s21[18], c21[18]);
	fa add2119(s20[20], a[19]&b[21], c21[18], s21[19], c21[19]);
	fa add2120(s20[21], a[20]&b[21], c21[19], s21[20], c21[20]);
	fa add2121(s20[22], a[21]&b[21], c21[20], s21[21], c21[21]);
	fa add2122(s20[23], a[22]&b[21], c21[21], s21[22], c21[22]);
	fa add2123(s20[24], a[23]&b[21], c21[22], s21[23], c21[23]);
	fa add2124(s20[25], a[24]&b[21], c21[23], s21[24], c21[24]);
	fa add2125(s20[26], a[25]&b[21], c21[24], s21[25], c21[25]);
	fa add2126(s20[27], a[26]&b[21], c21[25], s21[26], c21[26]);
	fa add2127(s20[28], a[27]&b[21], c21[26], s21[27], c21[27]);
	fa add2128(s20[29], a[28]&b[21], c21[27], s21[28], c21[28]);
	fa add2129(s20[30], a[29]&b[21], c21[28], s21[29], c21[29]);
	fa add2130(s20[31], a[30]&b[21], c21[29], s21[30], c21[30]);
	fa add2131(0, a[31]&b[21], c21[30], s21[31], c21[31]);
		
	
	wire [width-1:0] c22, s22;

	fa add2200(s21[1], a[0]&b[22], 0, prod[22], c22[0]);
	fa add2201(s21[2], a[1]&b[22], c22[0], s22[1], c22[1]);
	fa add2202(s21[3], a[2]&b[22], c22[1], s22[2], c22[2]);
	fa add2203(s21[4], a[3]&b[22], c22[2], s22[3], c22[3]);
	fa add2204(s21[5], a[4]&b[22], c22[3], s22[4], c22[4]);
	fa add2205(s21[6], a[5]&b[22], c22[4], s22[5], c22[5]);
	fa add2206(s21[7], a[6]&b[22], c22[5], s22[6], c22[6]);
	fa add2207(s21[8], a[7]&b[22], c22[6], s22[7], c22[7]);
	fa add2208(s21[9], a[8]&b[22], c22[7], s22[8], c22[8]);
	fa add2209(s21[10], a[9]&b[22], c22[8], s22[9], c22[9]);
	fa add2210(s21[11], a[10]&b[22], c22[9], s22[10], c22[10]);
	fa add2211(s21[12], a[11]&b[22], c22[10], s22[11], c22[11]);
	fa add2212(s21[13], a[12]&b[22], c22[11], s22[12], c22[12]);
	fa add2213(s21[14], a[13]&b[22], c22[12], s22[13], c22[13]);
	fa add2214(s21[15], a[14]&b[22], c22[13], s22[14], c22[14]);
	fa add2215(s21[16], a[15]&b[22], c22[14], s22[15], c22[15]);
	fa add2216(s21[17], a[16]&b[22], c22[15], s22[16], c22[16]);
	fa add2217(s21[18], a[17]&b[22], c22[16], s22[17], c22[17]);
	fa add2218(s21[19], a[18]&b[22], c22[17], s22[18], c22[18]);
	fa add2219(s21[20], a[19]&b[22], c22[18], s22[19], c22[19]);
	fa add2220(s21[21], a[20]&b[22], c22[19], s22[20], c22[20]);
	fa add2221(s21[22], a[21]&b[22], c22[20], s22[21], c22[21]);
	fa add2222(s21[23], a[22]&b[22], c22[21], s22[22], c22[22]);
	fa add2223(s21[24], a[23]&b[22], c22[22], s22[23], c22[23]);
	fa add2224(s21[25], a[24]&b[22], c22[23], s22[24], c22[24]);
	fa add2225(s21[26], a[25]&b[22], c22[24], s22[25], c22[25]);
	fa add2226(s21[27], a[26]&b[22], c22[25], s22[26], c22[26]);
	fa add2227(s21[28], a[27]&b[22], c22[26], s22[27], c22[27]);
	fa add2228(s21[29], a[28]&b[22], c22[27], s22[28], c22[28]);
	fa add2229(s21[30], a[29]&b[22], c22[28], s22[29], c22[29]);
	fa add2230(s21[31], a[30]&b[22], c22[29], s22[30], c22[30]);
	fa add2231(0, a[31]&b[22], c22[30], s22[31], c22[31]);
		
	
	wire [width-1:0] c23, s23;

	fa add2300(s22[1], a[0]&b[23], 0, prod[23], c23[0]);
	fa add2301(s22[2], a[1]&b[23], c23[0], s23[1], c23[1]);
	fa add2302(s22[3], a[2]&b[23], c23[1], s23[2], c23[2]);
	fa add2303(s22[4], a[3]&b[23], c23[2], s23[3], c23[3]);
	fa add2304(s22[5], a[4]&b[23], c23[3], s23[4], c23[4]);
	fa add2305(s22[6], a[5]&b[23], c23[4], s23[5], c23[5]);
	fa add2306(s22[7], a[6]&b[23], c23[5], s23[6], c23[6]);
	fa add2307(s22[8], a[7]&b[23], c23[6], s23[7], c23[7]);
	fa add2308(s22[9], a[8]&b[23], c23[7], s23[8], c23[8]);
	fa add2309(s22[10], a[9]&b[23], c23[8], s23[9], c23[9]);
	fa add2310(s22[11], a[10]&b[23], c23[9], s23[10], c23[10]);
	fa add2311(s22[12], a[11]&b[23], c23[10], s23[11], c23[11]);
	fa add2312(s22[13], a[12]&b[23], c23[11], s23[12], c23[12]);
	fa add2313(s22[14], a[13]&b[23], c23[12], s23[13], c23[13]);
	fa add2314(s22[15], a[14]&b[23], c23[13], s23[14], c23[14]);
	fa add2315(s22[16], a[15]&b[23], c23[14], s23[15], c23[15]);
	fa add2316(s22[17], a[16]&b[23], c23[15], s23[16], c23[16]);
	fa add2317(s22[18], a[17]&b[23], c23[16], s23[17], c23[17]);
	fa add2318(s22[19], a[18]&b[23], c23[17], s23[18], c23[18]);
	fa add2319(s22[20], a[19]&b[23], c23[18], s23[19], c23[19]);
	fa add2320(s22[21], a[20]&b[23], c23[19], s23[20], c23[20]);
	fa add2321(s22[22], a[21]&b[23], c23[20], s23[21], c23[21]);
	fa add2322(s22[23], a[22]&b[23], c23[21], s23[22], c23[22]);
	fa add2323(s22[24], a[23]&b[23], c23[22], s23[23], c23[23]);
	fa add2324(s22[25], a[24]&b[23], c23[23], s23[24], c23[24]);
	fa add2325(s22[26], a[25]&b[23], c23[24], s23[25], c23[25]);
	fa add2326(s22[27], a[26]&b[23], c23[25], s23[26], c23[26]);
	fa add2327(s22[28], a[27]&b[23], c23[26], s23[27], c23[27]);
	fa add2328(s22[29], a[28]&b[23], c23[27], s23[28], c23[28]);
	fa add2329(s22[30], a[29]&b[23], c23[28], s23[29], c23[29]);
	fa add2330(s22[31], a[30]&b[23], c23[29], s23[30], c23[30]);
	fa add2331(0, a[31]&b[23], c23[30], s23[31], c23[31]);
		
	
	wire [width-1:0] c24, s24;

	fa add2400(s23[1], a[0]&b[24], 0, prod[24], c24[0]);
	fa add2401(s23[2], a[1]&b[24], c24[0], s24[1], c24[1]);
	fa add2402(s23[3], a[2]&b[24], c24[1], s24[2], c24[2]);
	fa add2403(s23[4], a[3]&b[24], c24[2], s24[3], c24[3]);
	fa add2404(s23[5], a[4]&b[24], c24[3], s24[4], c24[4]);
	fa add2405(s23[6], a[5]&b[24], c24[4], s24[5], c24[5]);
	fa add2406(s23[7], a[6]&b[24], c24[5], s24[6], c24[6]);
	fa add2407(s23[8], a[7]&b[24], c24[6], s24[7], c24[7]);
	fa add2408(s23[9], a[8]&b[24], c24[7], s24[8], c24[8]);
	fa add2409(s23[10], a[9]&b[24], c24[8], s24[9], c24[9]);
	fa add2410(s23[11], a[10]&b[24], c24[9], s24[10], c24[10]);
	fa add2411(s23[12], a[11]&b[24], c24[10], s24[11], c24[11]);
	fa add2412(s23[13], a[12]&b[24], c24[11], s24[12], c24[12]);
	fa add2413(s23[14], a[13]&b[24], c24[12], s24[13], c24[13]);
	fa add2414(s23[15], a[14]&b[24], c24[13], s24[14], c24[14]);
	fa add2415(s23[16], a[15]&b[24], c24[14], s24[15], c24[15]);
	fa add2416(s23[17], a[16]&b[24], c24[15], s24[16], c24[16]);
	fa add2417(s23[18], a[17]&b[24], c24[16], s24[17], c24[17]);
	fa add2418(s23[19], a[18]&b[24], c24[17], s24[18], c24[18]);
	fa add2419(s23[20], a[19]&b[24], c24[18], s24[19], c24[19]);
	fa add2420(s23[21], a[20]&b[24], c24[19], s24[20], c24[20]);
	fa add2421(s23[22], a[21]&b[24], c24[20], s24[21], c24[21]);
	fa add2422(s23[23], a[22]&b[24], c24[21], s24[22], c24[22]);
	fa add2423(s23[24], a[23]&b[24], c24[22], s24[23], c24[23]);
	fa add2424(s23[25], a[24]&b[24], c24[23], s24[24], c24[24]);
	fa add2425(s23[26], a[25]&b[24], c24[24], s24[25], c24[25]);
	fa add2426(s23[27], a[26]&b[24], c24[25], s24[26], c24[26]);
	fa add2427(s23[28], a[27]&b[24], c24[26], s24[27], c24[27]);
	fa add2428(s23[29], a[28]&b[24], c24[27], s24[28], c24[28]);
	fa add2429(s23[30], a[29]&b[24], c24[28], s24[29], c24[29]);
	fa add2430(s23[31], a[30]&b[24], c24[29], s24[30], c24[30]);
	fa add2431(0, a[31]&b[24], c24[30], s24[31], c24[31]);
			
	
	wire [width-1:0] c25, s25;

	fa add2500(s24[1], a[0]&b[25], 0, prod[25], c25[0]);
	fa add2501(s24[2], a[1]&b[25], c25[0], s25[1], c25[1]);
	fa add2502(s24[3], a[2]&b[25], c25[1], s25[2], c25[2]);
	fa add2503(s24[4], a[3]&b[25], c25[2], s25[3], c25[3]);
	fa add2504(s24[5], a[4]&b[25], c25[3], s25[4], c25[4]);
	fa add2505(s24[6], a[5]&b[25], c25[4], s25[5], c25[5]);
	fa add2506(s24[7], a[6]&b[25], c25[5], s25[6], c25[6]);
	fa add2507(s24[8], a[7]&b[25], c25[6], s25[7], c25[7]);
	fa add2508(s24[9], a[8]&b[25], c25[7], s25[8], c25[8]);
	fa add2509(s24[10], a[9]&b[25], c25[8], s25[9], c25[9]);
	fa add2510(s24[11], a[10]&b[25], c25[9], s25[10], c25[10]);
	fa add2511(s24[12], a[11]&b[25], c25[10], s25[11], c25[11]);
	fa add2512(s24[13], a[12]&b[25], c25[11], s25[12], c25[12]);
	fa add2513(s24[14], a[13]&b[25], c25[12], s25[13], c25[13]);
	fa add2514(s24[15], a[14]&b[25], c25[13], s25[14], c25[14]);
	fa add2515(s24[16], a[15]&b[25], c25[14], s25[15], c25[15]);
	fa add2516(s24[17], a[16]&b[25], c25[15], s25[16], c25[16]);
	fa add2517(s24[18], a[17]&b[25], c25[16], s25[17], c25[17]);
	fa add2518(s24[19], a[18]&b[25], c25[17], s25[18], c25[18]);
	fa add2519(s24[20], a[19]&b[25], c25[18], s25[19], c25[19]);
	fa add2520(s24[21], a[20]&b[25], c25[19], s25[20], c25[20]);
	fa add2521(s24[22], a[21]&b[25], c25[20], s25[21], c25[21]);
	fa add2522(s24[23], a[22]&b[25], c25[21], s25[22], c25[22]);
	fa add2523(s24[24], a[23]&b[25], c25[22], s25[23], c25[23]);
	fa add2524(s24[25], a[24]&b[25], c25[23], s25[24], c25[24]);
	fa add2525(s24[26], a[25]&b[25], c25[24], s25[25], c25[25]);
	fa add2526(s24[27], a[26]&b[25], c25[25], s25[26], c25[26]);
	fa add2527(s24[28], a[27]&b[25], c25[26], s25[27], c25[27]);
	fa add2528(s24[29], a[28]&b[25], c25[27], s25[28], c25[28]);
	fa add2529(s24[30], a[29]&b[25], c25[28], s25[29], c25[29]);
	fa add2530(s24[31], a[30]&b[25], c25[29], s25[30], c25[30]);
	fa add2531(0, a[31]&b[25], c25[30], s25[31], c25[31]);
			
	
	wire [width-1:0] c26, s26;

	fa add2600(s25[1], a[0]&b[26], 0, prod[26], c26[0]);
	fa add2601(s25[2], a[1]&b[26], c26[0], s26[1], c26[1]);
	fa add2602(s25[3], a[2]&b[26], c26[1], s26[2], c26[2]);
	fa add2603(s25[4], a[3]&b[26], c26[2], s26[3], c26[3]);
	fa add2604(s25[5], a[4]&b[26], c26[3], s26[4], c26[4]);
	fa add2605(s25[6], a[5]&b[26], c26[4], s26[5], c26[5]);
	fa add2606(s25[7], a[6]&b[26], c26[5], s26[6], c26[6]);
	fa add2607(s25[8], a[7]&b[26], c26[6], s26[7], c26[7]);
	fa add2608(s25[9], a[8]&b[26], c26[7], s26[8], c26[8]);
	fa add2609(s25[10], a[9]&b[26], c26[8], s26[9], c26[9]);
	fa add2610(s25[11], a[10]&b[26], c26[9], s26[10], c26[10]);
	fa add2611(s25[12], a[11]&b[26], c26[10], s26[11], c26[11]);
	fa add2612(s25[13], a[12]&b[26], c26[11], s26[12], c26[12]);
	fa add2613(s25[14], a[13]&b[26], c26[12], s26[13], c26[13]);
	fa add2614(s25[15], a[14]&b[26], c26[13], s26[14], c26[14]);
	fa add2615(s25[16], a[15]&b[26], c26[14], s26[15], c26[15]);
	fa add2616(s25[17], a[16]&b[26], c26[15], s26[16], c26[16]);
	fa add2617(s25[18], a[17]&b[26], c26[16], s26[17], c26[17]);
	fa add2618(s25[19], a[18]&b[26], c26[17], s26[18], c26[18]);
	fa add2619(s25[20], a[19]&b[26], c26[18], s26[19], c26[19]);
	fa add2620(s25[21], a[20]&b[26], c26[19], s26[20], c26[20]);
	fa add2621(s25[22], a[21]&b[26], c26[20], s26[21], c26[21]);
	fa add2622(s25[23], a[22]&b[26], c26[21], s26[22], c26[22]);
	fa add2623(s25[24], a[23]&b[26], c26[22], s26[23], c26[23]);
	fa add2624(s25[25], a[24]&b[26], c26[23], s26[24], c26[24]);
	fa add2625(s25[26], a[25]&b[26], c26[24], s26[25], c26[25]);
	fa add2626(s25[27], a[26]&b[26], c26[25], s26[26], c26[26]);
	fa add2627(s25[28], a[27]&b[26], c26[26], s26[27], c26[27]);
	fa add2628(s25[29], a[28]&b[26], c26[27], s26[28], c26[28]);
	fa add2629(s25[30], a[29]&b[26], c26[28], s26[29], c26[29]);
	fa add2630(s25[31], a[30]&b[26], c26[29], s26[30], c26[30]);
	fa add2631(0, a[31]&b[26], c26[30], s26[31], c26[31]);
			
	
	wire [width-1:0] c27, s27;

	fa add2700(s26[1], a[0]&b[27], 0, prod[27], c27[0]);
	fa add2701(s26[2], a[1]&b[27], c27[0], s27[1], c27[1]);
	fa add2702(s26[3], a[2]&b[27], c27[1], s27[2], c27[2]);
	fa add2703(s26[4], a[3]&b[27], c27[2], s27[3], c27[3]);
	fa add2704(s26[5], a[4]&b[27], c27[3], s27[4], c27[4]);
	fa add2705(s26[6], a[5]&b[27], c27[4], s27[5], c27[5]);
	fa add2706(s26[7], a[6]&b[27], c27[5], s27[6], c27[6]);
	fa add2707(s26[8], a[7]&b[27], c27[6], s27[7], c27[7]);
	fa add2708(s26[9], a[8]&b[27], c27[7], s27[8], c27[8]);
	fa add2709(s26[10], a[9]&b[27], c27[8], s27[9], c27[9]);
	fa add2710(s26[11], a[10]&b[27], c27[9], s27[10], c27[10]);
	fa add2711(s26[12], a[11]&b[27], c27[10], s27[11], c27[11]);
	fa add2712(s26[13], a[12]&b[27], c27[11], s27[12], c27[12]);
	fa add2713(s26[14], a[13]&b[27], c27[12], s27[13], c27[13]);
	fa add2714(s26[15], a[14]&b[27], c27[13], s27[14], c27[14]);
	fa add2715(s26[16], a[15]&b[27], c27[14], s27[15], c27[15]);
	fa add2716(s26[17], a[16]&b[27], c27[15], s27[16], c27[16]);
	fa add2717(s26[18], a[17]&b[27], c27[16], s27[17], c27[17]);
	fa add2718(s26[19], a[18]&b[27], c27[17], s27[18], c27[18]);
	fa add2719(s26[20], a[19]&b[27], c27[18], s27[19], c27[19]);
	fa add2720(s26[21], a[20]&b[27], c27[19], s27[20], c27[20]);
	fa add2721(s26[22], a[21]&b[27], c27[20], s27[21], c27[21]);
	fa add2722(s26[23], a[22]&b[27], c27[21], s27[22], c27[22]);
	fa add2723(s26[24], a[23]&b[27], c27[22], s27[23], c27[23]);
	fa add2724(s26[25], a[24]&b[27], c27[23], s27[24], c27[24]);
	fa add2725(s26[26], a[25]&b[27], c27[24], s27[25], c27[25]);
	fa add2726(s26[27], a[26]&b[27], c27[25], s27[26], c27[26]);
	fa add2727(s26[28], a[27]&b[27], c27[26], s27[27], c27[27]);
	fa add2728(s26[29], a[28]&b[27], c27[27], s27[28], c27[28]);
	fa add2729(s26[30], a[29]&b[27], c27[28], s27[29], c27[29]);
	fa add2730(s26[31], a[30]&b[27], c27[29], s27[30], c27[30]);
	fa add2731(0, a[31]&b[27], c27[30], s27[31], c27[31]);
			
	
	wire [width-1:0] c28, s28;

	fa add2800(s27[1], a[0]&b[28], 0, prod[28], c28[0]);
	fa add2801(s27[2], a[1]&b[28], c28[0], s28[1], c28[1]);
	fa add2802(s27[3], a[2]&b[28], c28[1], s28[2], c28[2]);
	fa add2803(s27[4], a[3]&b[28], c28[2], s28[3], c28[3]);
	fa add2804(s27[5], a[4]&b[28], c28[3], s28[4], c28[4]);
	fa add2805(s27[6], a[5]&b[28], c28[4], s28[5], c28[5]);
	fa add2806(s27[7], a[6]&b[28], c28[5], s28[6], c28[6]);
	fa add2807(s27[8], a[7]&b[28], c28[6], s28[7], c28[7]);
	fa add2808(s27[9], a[8]&b[28], c28[7], s28[8], c28[8]);
	fa add2809(s27[10], a[9]&b[28], c28[8], s28[9], c28[9]);
	fa add2810(s27[11], a[10]&b[28], c28[9], s28[10], c28[10]);
	fa add2811(s27[12], a[11]&b[28], c28[10], s28[11], c28[11]);
	fa add2812(s27[13], a[12]&b[28], c28[11], s28[12], c28[12]);
	fa add2813(s27[14], a[13]&b[28], c28[12], s28[13], c28[13]);
	fa add2814(s27[15], a[14]&b[28], c28[13], s28[14], c28[14]);
	fa add2815(s27[16], a[15]&b[28], c28[14], s28[15], c28[15]);
	fa add2816(s27[17], a[16]&b[28], c28[15], s28[16], c28[16]);
	fa add2817(s27[18], a[17]&b[28], c28[16], s28[17], c28[17]);
	fa add2818(s27[19], a[18]&b[28], c28[17], s28[18], c28[18]);
	fa add2819(s27[20], a[19]&b[28], c28[18], s28[19], c28[19]);
	fa add2820(s27[21], a[20]&b[28], c28[19], s28[20], c28[20]);
	fa add2821(s27[22], a[21]&b[28], c28[20], s28[21], c28[21]);
	fa add2822(s27[23], a[22]&b[28], c28[21], s28[22], c28[22]);
	fa add2823(s27[24], a[23]&b[28], c28[22], s28[23], c28[23]);
	fa add2824(s27[25], a[24]&b[28], c28[23], s28[24], c28[24]);
	fa add2825(s27[26], a[25]&b[28], c28[24], s28[25], c28[25]);
	fa add2826(s27[27], a[26]&b[28], c28[25], s28[26], c28[26]);
	fa add2827(s27[28], a[27]&b[28], c28[26], s28[27], c28[27]);
	fa add2828(s27[29], a[28]&b[28], c28[27], s28[28], c28[28]);
	fa add2829(s27[30], a[29]&b[28], c28[28], s28[29], c28[29]);
	fa add2830(s27[31], a[30]&b[28], c28[29], s28[30], c28[30]);
	fa add2831(0, a[31]&b[28], c28[30], s28[31], c28[31]);
			
	
	wire [width-1:0] c29, s29;

	fa add2900(s28[1], a[0]&b[29], 0, prod[29], c29[0]);
	fa add2901(s28[2], a[1]&b[29], c29[0], s29[1], c29[1]);
	fa add2902(s28[3], a[2]&b[29], c29[1], s29[2], c29[2]);
	fa add2903(s28[4], a[3]&b[29], c29[2], s29[3], c29[3]);
	fa add2904(s28[5], a[4]&b[29], c29[3], s29[4], c29[4]);
	fa add2905(s28[6], a[5]&b[29], c29[4], s29[5], c29[5]);
	fa add2906(s28[7], a[6]&b[29], c29[5], s29[6], c29[6]);
	fa add2907(s28[8], a[7]&b[29], c29[6], s29[7], c29[7]);
	fa add2908(s28[9], a[8]&b[29], c29[7], s29[8], c29[8]);
	fa add2909(s28[10], a[9]&b[29], c29[8], s29[9], c29[9]);
	fa add2910(s28[11], a[10]&b[29], c29[9], s29[10], c29[10]);
	fa add2911(s28[12], a[11]&b[29], c29[10], s29[11], c29[11]);
	fa add2912(s28[13], a[12]&b[29], c29[11], s29[12], c29[12]);
	fa add2913(s28[14], a[13]&b[29], c29[12], s29[13], c29[13]);
	fa add2914(s28[15], a[14]&b[29], c29[13], s29[14], c29[14]);
	fa add2915(s28[16], a[15]&b[29], c29[14], s29[15], c29[15]);
	fa add2916(s28[17], a[16]&b[29], c29[15], s29[16], c29[16]);
	fa add2917(s28[18], a[17]&b[29], c29[16], s29[17], c29[17]);
	fa add2918(s28[19], a[18]&b[29], c29[17], s29[18], c29[18]);
	fa add2919(s28[20], a[19]&b[29], c29[18], s29[19], c29[19]);
	fa add2920(s28[21], a[20]&b[29], c29[19], s29[20], c29[20]);
	fa add2921(s28[22], a[21]&b[29], c29[20], s29[21], c29[21]);
	fa add2922(s28[23], a[22]&b[29], c29[21], s29[22], c29[22]);
	fa add2923(s28[24], a[23]&b[29], c29[22], s29[23], c29[23]);
	fa add2924(s28[25], a[24]&b[29], c29[23], s29[24], c29[24]);
	fa add2925(s28[26], a[25]&b[29], c29[24], s29[25], c29[25]);
	fa add2926(s28[27], a[26]&b[29], c29[25], s29[26], c29[26]);
	fa add2927(s28[28], a[27]&b[29], c29[26], s29[27], c29[27]);
	fa add2928(s28[29], a[28]&b[29], c29[27], s29[28], c29[28]);
	fa add2929(s28[30], a[29]&b[29], c29[28], s29[29], c29[29]);
	fa add2930(s28[31], a[30]&b[29], c29[29], s29[30], c29[30]);
	fa add2931(0, a[31]&b[29], c29[30], s29[31], c29[31]);
			
	
	wire [width-1:0] c30, s30;

	fa add3000(s29[1], a[0]&b[30], 0, prod[30], c30[0]);
	fa add3001(s29[2], a[1]&b[30], c30[0], s30[1], c30[1]);
	fa add3002(s29[3], a[2]&b[30], c30[1], s30[2], c30[2]);
	fa add3003(s29[4], a[3]&b[30], c30[2], s30[3], c30[3]);
	fa add3004(s29[5], a[4]&b[30], c30[3], s30[4], c30[4]);
	fa add3005(s29[6], a[5]&b[30], c30[4], s30[5], c30[5]);
	fa add3006(s29[7], a[6]&b[30], c30[5], s30[6], c30[6]);
	fa add3007(s29[8], a[7]&b[30], c30[6], s30[7], c30[7]);
	fa add3008(s29[9], a[8]&b[30], c30[7], s30[8], c30[8]);
	fa add3009(s29[10], a[9]&b[30], c30[8], s30[9], c30[9]);
	fa add3010(s29[11], a[10]&b[30], c30[9], s30[10], c30[10]);
	fa add3011(s29[12], a[11]&b[30], c30[10], s30[11], c30[11]);
	fa add3012(s29[13], a[12]&b[30], c30[11], s30[12], c30[12]);
	fa add3013(s29[14], a[13]&b[30], c30[12], s30[13], c30[13]);
	fa add3014(s29[15], a[14]&b[30], c30[13], s30[14], c30[14]);
	fa add3015(s29[16], a[15]&b[30], c30[14], s30[15], c30[15]);
	fa add3016(s29[17], a[16]&b[30], c30[15], s30[16], c30[16]);
	fa add3017(s29[18], a[17]&b[30], c30[16], s30[17], c30[17]);
	fa add3018(s29[19], a[18]&b[30], c30[17], s30[18], c30[18]);
	fa add3019(s29[20], a[19]&b[30], c30[18], s30[19], c30[19]);
	fa add3020(s29[21], a[20]&b[30], c30[19], s30[20], c30[20]);
	fa add3021(s29[22], a[21]&b[30], c30[20], s30[21], c30[21]);
	fa add3022(s29[23], a[22]&b[30], c30[21], s30[22], c30[22]);
	fa add3023(s29[24], a[23]&b[30], c30[22], s30[23], c30[23]);
	fa add3024(s29[25], a[24]&b[30], c30[23], s30[24], c30[24]);
	fa add3025(s29[26], a[25]&b[30], c30[24], s30[25], c30[25]);
	fa add3026(s29[27], a[26]&b[30], c30[25], s30[26], c30[26]);
	fa add3027(s29[28], a[27]&b[30], c30[26], s30[27], c30[27]);
	fa add3028(s29[29], a[28]&b[30], c30[27], s30[28], c30[28]);
	fa add3029(s29[30], a[29]&b[30], c30[28], s30[29], c30[29]);
	fa add3030(s29[31], a[30]&b[30], c30[29], s30[30], c30[30]);
	fa add3031(0, a[31]&b[30], c30[30], s30[31], c30[31]);
			
	
	wire [width-1:0] c31, s31;

	fa add3100(s30[1], a[0]&b[31], 0, prod[31], c31[0]);
	fa add3101(s30[2], a[1]&b[31], c31[0], s31[1], c31[1]);
	fa add3102(s30[3], a[2]&b[31], c31[1], s31[2], c31[2]);
	fa add3103(s30[4], a[3]&b[31], c31[2], s31[3], c31[3]);
	fa add3104(s30[5], a[4]&b[31], c31[3], s31[4], c31[4]);
	fa add3105(s30[6], a[5]&b[31], c31[4], s31[5], c31[5]);
	fa add3106(s30[7], a[6]&b[31], c31[5], s31[6], c31[6]);
	fa add3107(s30[8], a[7]&b[31], c31[6], s31[7], c31[7]);
	fa add3108(s30[9], a[8]&b[31], c31[7], s31[8], c31[8]);
	fa add3109(s30[10], a[9]&b[31], c31[8], s31[9], c31[9]);
	fa add3110(s30[11], a[10]&b[31], c31[9], s31[10], c31[10]);
	fa add3111(s30[12], a[11]&b[31], c31[10], s31[11], c31[11]);
	fa add3112(s30[13], a[12]&b[31], c31[11], s31[12], c31[12]);
	fa add3113(s30[14], a[13]&b[31], c31[12], s31[13], c31[13]);
	fa add3114(s30[15], a[14]&b[31], c31[13], s31[14], c31[14]);
	fa add3115(s30[16], a[15]&b[31], c31[14], s31[15], c31[15]);
	fa add3116(s30[17], a[16]&b[31], c31[15], s31[16], c31[16]);
	fa add3117(s30[18], a[17]&b[31], c31[16], s31[17], c31[17]);
	fa add3118(s30[19], a[18]&b[31], c31[17], s31[18], c31[18]);
	fa add3119(s30[20], a[19]&b[31], c31[18], s31[19], c31[19]);
	fa add3120(s30[21], a[20]&b[31], c31[19], s31[20], c31[20]);
	fa add3121(s30[22], a[21]&b[31], c31[20], s31[21], c31[21]);
	fa add3122(s30[23], a[22]&b[31], c31[21], s31[22], c31[22]);
	fa add3123(s30[24], a[23]&b[31], c31[22], s31[23], c31[23]);
	fa add3124(s30[25], a[24]&b[31], c31[23], s31[24], c31[24]);
	fa add3125(s30[26], a[25]&b[31], c31[24], s31[25], c31[25]);
	fa add3126(s30[27], a[26]&b[31], c31[25], s31[26], c31[26]);
	fa add3127(s30[28], a[27]&b[31], c31[26], s31[27], c31[27]);
	fa add3128(s30[29], a[28]&b[31], c31[27], s31[28], c31[28]);
	fa add3129(s30[30], a[29]&b[31], c31[28], s31[29], c31[29]);
	fa add3130(s30[31], a[30]&b[31], c31[29], s31[30], c31[30]);
	fa add3131(0, a[31]&b[31], c31[30], s31[31], c31[31]);

endmodule
