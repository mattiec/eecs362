module 32b_slt(a,b,c);
	parameter width = 32;

	input [0:width-1] a,b;
	output c;

endmodule
